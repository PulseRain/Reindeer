module single_port_ram_sim_high #(parameter ADDR_WIDTH, DATA_WIDTH ) (
    input  wire [ADDR_WIDTH - 1 : 0]         addr,
    input  wire [DATA_WIDTH - 1 : 0]         din,
    input  wire [DATA_WIDTH / 8 - 1 : 0]     write_en,
    input  wire                              clk,
    output reg [DATA_WIDTH - 1 : 0]          dout
);
    reg [DATA_WIDTH - 1 : 0] mem [(1<<ADDR_WIDTH)-1:0];
    genvar i;
    generate
        for (i = 0; i < (DATA_WIDTH / 8); i = i + 1) begin : gen_proc
            always @(posedge clk) begin
                if (write_en[i]) begin
                    mem[(addr)][8 * (i + 1) - 1 : 8 * i] <= din[8 * (i + 1) - 1 : 8 * i];
                end
            end
        end
    endgenerate
 
    always @(posedge clk) begin
        dout <= mem[addr];
    end
 
initial begin
//================================================================
//== Section  .note.gnu.build-id
//================================================================
    mem[0] <= 16'h0000; // 0x80000000
    mem[1] <= 16'h0000; // 0x80000004
    mem[2] <= 16'h0000; // 0x80000008
    mem[3] <= 16'h0055; // 0x8000000c
    mem[4] <= 16'h1bfa; // 0x80000010
    mem[5] <= 16'hf88e; // 0x80000014
    mem[6] <= 16'hd3f2; // 0x80000018
    mem[7] <= 16'h79b4; // 0x8000001c
    mem[8] <= 16'h9bc4; // 0x80000020
 
 
//================================================================
//== Section  .text.init
//================================================================
    mem[9] <= 16'h0000; // 0x80000024
    mem[10] <= 16'h0000; // 0x80000028
    mem[11] <= 16'h0000; // 0x8000002c
    mem[12] <= 16'h0000; // 0x80000030
    mem[13] <= 16'h0000; // 0x80000034
    mem[14] <= 16'h0000; // 0x80000038
    mem[15] <= 16'h0000; // 0x8000003c
    mem[16] <= 16'h0000; // 0x80000040
    mem[17] <= 16'h0000; // 0x80000044
    mem[18] <= 16'h0000; // 0x80000048
    mem[19] <= 16'h0000; // 0x8000004c
    mem[20] <= 16'h0000; // 0x80000050
    mem[21] <= 16'h0000; // 0x80000054
    mem[22] <= 16'h0000; // 0x80000058
    mem[23] <= 16'h0000; // 0x8000005c
    mem[24] <= 16'h0000; // 0x80000060
    mem[25] <= 16'h0000; // 0x80000064
    mem[26] <= 16'h0000; // 0x80000068
    mem[27] <= 16'h0000; // 0x8000006c
    mem[28] <= 16'h0000; // 0x80000070
    mem[29] <= 16'h0000; // 0x80000074
    mem[30] <= 16'h0000; // 0x80000078
    mem[31] <= 16'h0000; // 0x8000007c
    mem[32] <= 16'h0000; // 0x80000080
    mem[33] <= 16'h0000; // 0x80000084
    mem[34] <= 16'h0000; // 0x80000088
    mem[35] <= 16'h0000; // 0x8000008c
    mem[36] <= 16'h0000; // 0x80000090
    mem[37] <= 16'h0000; // 0x80000094
    mem[38] <= 16'h0000; // 0x80000098
    mem[39] <= 16'h0000; // 0x8000009c
    mem[40] <= 16'h0001; // 0x800000a0
    mem[41] <= 16'h3002; // 0x800000a4
    mem[42] <= 16'h0010; // 0x800000a8
    mem[43] <= 16'h01f2; // 0x800000ac
    mem[44] <= 16'h0002; // 0x800000b0
    mem[45] <= 16'h0010; // 0x800000b4
    mem[46] <= 16'h0000; // 0x800000b8
    mem[47] <= 16'hf4a2; // 0x800000bc
    mem[48] <= 16'hff5f; // 0x800000c0
    mem[49] <= 16'h0000; // 0x800000c4
    mem[50] <= 16'h0442; // 0x800000c8
    mem[51] <= 16'h3052; // 0x800000cc
    mem[52] <= 16'h0000; // 0x800000d0
    mem[53] <= 16'hbec1; // 0x800000d4
    mem[54] <= 16'h0000; // 0x800000d8
    mem[55] <= 16'hc472; // 0x800000dc
    mem[56] <= 16'hfc02; // 0x800000e0
    mem[57] <= 16'hf140; // 0x800000e4
    mem[58] <= 16'h0010; // 0x800000e8
    mem[59] <= 16'h00b5; // 0x800000ec
    mem[60] <= 16'h00c5; // 0x800000f0
    mem[61] <= 16'h00c2; // 0x800000f4
    mem[62] <= 16'h0015; // 0x800000f8
    mem[63] <= 16'h00c1; // 0x800000fc
    mem[64] <= 16'h0041; // 0x80000100
    mem[65] <= 16'h0d00; // 0x80000104
    mem[66] <= 16'hef01; // 0x80000108
    mem[67] <= 16'h0011; // 0x8000010c
    mem[68] <= 16'h0021; // 0x80000110
    mem[69] <= 16'h0031; // 0x80000114
    mem[70] <= 16'h0041; // 0x80000118
    mem[71] <= 16'h0051; // 0x8000011c
    mem[72] <= 16'h0061; // 0x80000120
    mem[73] <= 16'h0071; // 0x80000124
    mem[74] <= 16'h0281; // 0x80000128
    mem[75] <= 16'h0291; // 0x8000012c
    mem[76] <= 16'h02a1; // 0x80000130
    mem[77] <= 16'h02b1; // 0x80000134
    mem[78] <= 16'h02c1; // 0x80000138
    mem[79] <= 16'h02d1; // 0x8000013c
    mem[80] <= 16'h02e1; // 0x80000140
    mem[81] <= 16'h02f1; // 0x80000144
    mem[82] <= 16'h0501; // 0x80000148
    mem[83] <= 16'h0511; // 0x8000014c
    mem[84] <= 16'h0521; // 0x80000150
    mem[85] <= 16'h0531; // 0x80000154
    mem[86] <= 16'h0541; // 0x80000158
    mem[87] <= 16'h0551; // 0x8000015c
    mem[88] <= 16'h0561; // 0x80000160
    mem[89] <= 16'h0571; // 0x80000164
    mem[90] <= 16'h0781; // 0x80000168
    mem[91] <= 16'h0791; // 0x8000016c
    mem[92] <= 16'h07a1; // 0x80000170
    mem[93] <= 16'h07b1; // 0x80000174
    mem[94] <= 16'h07c1; // 0x80000178
    mem[95] <= 16'h07d1; // 0x8000017c
    mem[96] <= 16'h07e1; // 0x80000180
    mem[97] <= 16'h07f1; // 0x80000184
    mem[98] <= 16'h3420; // 0x80000188
    mem[99] <= 16'h3410; // 0x8000018c
    mem[100] <= 16'h0001; // 0x80000190
    mem[101] <= 16'h6e80; // 0x80000194
    mem[102] <= 16'h3415; // 0x80000198
    mem[103] <= 16'h0000; // 0x8000019c
    mem[104] <= 16'h8002; // 0x800001a0
    mem[105] <= 16'h3002; // 0x800001a4
    mem[106] <= 16'h0041; // 0x800001a8
    mem[107] <= 16'h0081; // 0x800001ac
    mem[108] <= 16'h00c1; // 0x800001b0
    mem[109] <= 16'h0101; // 0x800001b4
    mem[110] <= 16'h0141; // 0x800001b8
    mem[111] <= 16'h0181; // 0x800001bc
    mem[112] <= 16'h01c1; // 0x800001c0
    mem[113] <= 16'h0201; // 0x800001c4
    mem[114] <= 16'h0241; // 0x800001c8
    mem[115] <= 16'h0281; // 0x800001cc
    mem[116] <= 16'h02c1; // 0x800001d0
    mem[117] <= 16'h0301; // 0x800001d4
    mem[118] <= 16'h0341; // 0x800001d8
    mem[119] <= 16'h0381; // 0x800001dc
    mem[120] <= 16'h03c1; // 0x800001e0
    mem[121] <= 16'h0401; // 0x800001e4
    mem[122] <= 16'h0441; // 0x800001e8
    mem[123] <= 16'h0481; // 0x800001ec
    mem[124] <= 16'h04c1; // 0x800001f0
    mem[125] <= 16'h0501; // 0x800001f4
    mem[126] <= 16'h0541; // 0x800001f8
    mem[127] <= 16'h0581; // 0x800001fc
    mem[128] <= 16'h05c1; // 0x80000200
    mem[129] <= 16'h0601; // 0x80000204
    mem[130] <= 16'h0641; // 0x80000208
    mem[131] <= 16'h0681; // 0x8000020c
    mem[132] <= 16'h06c1; // 0x80000210
    mem[133] <= 16'h0701; // 0x80000214
    mem[134] <= 16'h0741; // 0x80000218
    mem[135] <= 16'h0781; // 0x8000021c
    mem[136] <= 16'h07c1; // 0x80000220
    mem[137] <= 16'h1101; // 0x80000224
    mem[138] <= 16'h3020; // 0x80000228
 
 
//================================================================
//== Section  .tohost
//================================================================
    mem[1024] <= 16'h0000; // 0x80001000
    mem[1025] <= 16'h0000; // 0x80001004
    mem[1026] <= 16'h0000; // 0x80001008
    mem[1027] <= 16'h0000; // 0x8000100c
    mem[1028] <= 16'h0000; // 0x80001010
    mem[1029] <= 16'h0000; // 0x80001014
    mem[1030] <= 16'h0000; // 0x80001018
    mem[1031] <= 16'h0000; // 0x8000101c
    mem[1032] <= 16'h0000; // 0x80001020
    mem[1033] <= 16'h0000; // 0x80001024
    mem[1034] <= 16'h0000; // 0x80001028
    mem[1035] <= 16'h0000; // 0x8000102c
    mem[1036] <= 16'h0000; // 0x80001030
    mem[1037] <= 16'h0000; // 0x80001034
    mem[1038] <= 16'h0000; // 0x80001038
    mem[1039] <= 16'h0000; // 0x8000103c
    mem[1040] <= 16'h0000; // 0x80001040
    mem[1041] <= 16'h0000; // 0x80001044
 
 
//================================================================
//== Section  .text
//================================================================
    mem[1042] <= 16'h0025; // 0x80001048
    mem[1043] <= 16'h00b5; // 0x8000104c
    mem[1044] <= 16'h00b6; // 0x80001050
    mem[1045] <= 16'h0000; // 0x80001054
    mem[1046] <= 16'hfe01; // 0x80001058
    mem[1047] <= 16'h0131; // 0x8000105c
    mem[1048] <= 16'h0056; // 0x80001060
    mem[1049] <= 16'h0091; // 0x80001064
    mem[1050] <= 16'h0029; // 0x80001068
    mem[1051] <= 16'h0011; // 0x8000106c
    mem[1052] <= 16'h0081; // 0x80001070
    mem[1053] <= 16'h0121; // 0x80001074
    mem[1054] <= 16'h0095; // 0x80001078
    mem[1055] <= 16'h0005; // 0x8000107c
    mem[1056] <= 16'h0734; // 0x80001080
    mem[1057] <= 16'h0006; // 0x80001084
    mem[1058] <= 16'h00d4; // 0x80001088
    mem[1059] <= 16'h00d4; // 0x8000108c
    mem[1060] <= 16'h0009; // 0x80001090
    mem[1061] <= 16'h0c80; // 0x80001094
    mem[1062] <= 16'h7890; // 0x80001098
    mem[1063] <= 16'h0029; // 0x8000109c
    mem[1064] <= 16'h0125; // 0x800010a0
    mem[1065] <= 16'h00f4; // 0x800010a4
    mem[1066] <= 16'h0107; // 0x800010a8
    mem[1067] <= 16'h0137; // 0x800010ac
    mem[1068] <= 16'h0137; // 0x800010b0
    mem[1069] <= 16'h0017; // 0x800010b4
    mem[1070] <= 16'h00e7; // 0x800010b8
    mem[1071] <= 16'h0004; // 0x800010bc
    mem[1072] <= 16'h00a4; // 0x800010c0
    mem[1073] <= 16'h01c1; // 0x800010c4
    mem[1074] <= 16'h0124; // 0x800010c8
    mem[1075] <= 16'h0000; // 0x800010cc
    mem[1076] <= 16'h0087; // 0x800010d0
    mem[1077] <= 16'h0050; // 0x800010d4
    mem[1078] <= 16'hfae4; // 0x800010d8
    mem[1079] <= 16'h0141; // 0x800010dc
    mem[1080] <= 16'h0181; // 0x800010e0
    mem[1081] <= 16'h0101; // 0x800010e4
    mem[1082] <= 16'h00c1; // 0x800010e8
    mem[1083] <= 16'h0000; // 0x800010ec
    mem[1084] <= 16'h40f2; // 0x800010f0
    mem[1085] <= 16'h0201; // 0x800010f4
    mem[1086] <= 16'h0000; // 0x800010f8
    mem[1087] <= 16'h0ff5; // 0x800010fc
    mem[1088] <= 16'h0ff5; // 0x80001100
    mem[1089] <= 16'h00b5; // 0x80001104
    mem[1090] <= 16'h0000; // 0x80001108
    mem[1091] <= 16'h0000; // 0x8000110c
    mem[1092] <= 16'h0000; // 0x80001110
    mem[1093] <= 16'h3ca2; // 0x80001114
    mem[1094] <= 16'h0010; // 0x80001118
    mem[1095] <= 16'h0000; // 0x8000111c
    mem[1096] <= 16'hff01; // 0x80001120
    mem[1097] <= 16'h0081; // 0x80001124
    mem[1098] <= 16'h0091; // 0x80001128
    mem[1099] <= 16'h0011; // 0x8000112c
    mem[1100] <= 16'h0005; // 0x80001130
    mem[1101] <= 16'h0005; // 0x80001134
    mem[1102] <= 16'h0034; // 0x80001138
    mem[1103] <= 16'h0024; // 0x8000113c
    mem[1104] <= 16'hfbdf; // 0x80001140
    mem[1105] <= 16'hfe05; // 0x80001144
    mem[1106] <= 16'h0004; // 0x80001148
    mem[1107] <= 16'h0004; // 0x8000114c
    mem[1108] <= 16'h5640; // 0x80001150
    mem[1109] <= 16'h02a0; // 0x80001154
    mem[1110] <= 16'h00c1; // 0x80001158
    mem[1111] <= 16'h00a0; // 0x8000115c
    mem[1112] <= 16'h0010; // 0x80001160
    mem[1113] <= 16'h0081; // 0x80001164
    mem[1114] <= 16'h0041; // 0x80001168
    mem[1115] <= 16'h0000; // 0x8000116c
    mem[1116] <= 16'h38f2; // 0x80001170
    mem[1117] <= 16'h0101; // 0x80001174
    mem[1118] <= 16'h0000; // 0x80001178
    mem[1119] <= 16'h00c1; // 0x8000117c
    mem[1120] <= 16'h0000; // 0x80001180
    mem[1121] <= 16'h0081; // 0x80001184
    mem[1122] <= 16'h0041; // 0x80001188
    mem[1123] <= 16'h0101; // 0x8000118c
    mem[1124] <= 16'h0000; // 0x80001190
    mem[1125] <= 16'hffe5; // 0x80001194
    mem[1126] <= 16'h0015; // 0x80001198
    mem[1127] <= 16'h0000; // 0x8000119c
    mem[1128] <= 16'hff01; // 0x800011a0
    mem[1129] <= 16'h0081; // 0x800011a4
    mem[1130] <= 16'h0091; // 0x800011a8
    mem[1131] <= 16'h0011; // 0x800011ac
    mem[1132] <= 16'h0005; // 0x800011b0
    mem[1133] <= 16'h0005; // 0x800011b4
    mem[1134] <= 16'hfddf; // 0x800011b8
    mem[1135] <= 16'h0205; // 0x800011bc
    mem[1136] <= 16'h0084; // 0x800011c0
    mem[1137] <= 16'h0010; // 0x800011c4
    mem[1138] <= 16'h04f4; // 0x800011c8
    mem[1139] <= 16'h0404; // 0x800011cc
    mem[1140] <= 16'h0020; // 0x800011d0
    mem[1141] <= 16'h04e4; // 0x800011d4
    mem[1142] <= 16'h0040; // 0x800011d8
    mem[1143] <= 16'h00f4; // 0x800011dc
    mem[1144] <= 16'h00e4; // 0x800011e0
    mem[1145] <= 16'h00c1; // 0x800011e4
    mem[1146] <= 16'h0081; // 0x800011e8
    mem[1147] <= 16'h0041; // 0x800011ec
    mem[1148] <= 16'h0101; // 0x800011f0
    mem[1149] <= 16'h0000; // 0x800011f4
    mem[1150] <= 16'h0030; // 0x800011f8
    mem[1151] <= 16'h00f4; // 0x800011fc
    mem[1152] <= 16'h0010; // 0x80001200
    mem[1153] <= 16'hfcf4; // 0x80001204
    mem[1154] <= 16'h0000; // 0x80001208
    mem[1155] <= 16'h2e47; // 0x8000120c
    mem[1156] <= 16'h0640; // 0x80001210
    mem[1157] <= 16'h02e7; // 0x80001214
    mem[1158] <= 16'h00c1; // 0x80001218
    mem[1159] <= 16'h0004; // 0x8000121c
    mem[1160] <= 16'h0081; // 0x80001220
    mem[1161] <= 16'h0041; // 0x80001224
    mem[1162] <= 16'h0101; // 0x80001228
    mem[1163] <= 16'h0000; // 0x8000122c
    mem[1164] <= 16'h00c1; // 0x80001230
    mem[1165] <= 16'h00f4; // 0x80001234
    mem[1166] <= 16'h0081; // 0x80001238
    mem[1167] <= 16'h0041; // 0x8000123c
    mem[1168] <= 16'h0101; // 0x80001240
    mem[1169] <= 16'h0000; // 0x80001244
    mem[1170] <= 16'h00c1; // 0x80001248
    mem[1171] <= 16'h0030; // 0x8000124c
    mem[1172] <= 16'h00f4; // 0x80001250
    mem[1173] <= 16'h0081; // 0x80001254
    mem[1174] <= 16'h0041; // 0x80001258
    mem[1175] <= 16'h0101; // 0x8000125c
    mem[1176] <= 16'h0000; // 0x80001260
    mem[1177] <= 16'h0000; // 0x80001264
    mem[1178] <= 16'h2817; // 0x80001268
    mem[1179] <= 16'h0410; // 0x8000126c
    mem[1180] <= 16'h00f7; // 0x80001270
    mem[1181] <= 16'h0000; // 0x80001274
    mem[1182] <= 16'h0005; // 0x80001278
    mem[1183] <= 16'h0000; // 0x8000127c
    mem[1184] <= 16'h2707; // 0x80001280
    mem[1185] <= 16'h0097; // 0x80001284
    mem[1186] <= 16'h40e7; // 0x80001288
    mem[1187] <= 16'h00f5; // 0x8000128c
    mem[1188] <= 16'h0000; // 0x80001290
    mem[1189] <= 16'h0000; // 0x80001294
    mem[1190] <= 16'h2606; // 0x80001298
    mem[1191] <= 16'h0006; // 0x8000129c
    mem[1192] <= 16'h0006; // 0x800012a0
    mem[1193] <= 16'h00f5; // 0x800012a4
    mem[1194] <= 16'h0000; // 0x800012a8
    mem[1195] <= 16'h24c6; // 0x800012ac
    mem[1196] <= 16'h00c6; // 0x800012b0
    mem[1197] <= 16'h0000; // 0x800012b4
    mem[1198] <= 16'h2385; // 0x800012b8
    mem[1199] <= 16'h00a0; // 0x800012bc
    mem[1200] <= 16'hd89f; // 0x800012c0
    mem[1201] <= 16'h0000; // 0x800012c4
    mem[1202] <= 16'h2307; // 0x800012c8
    mem[1203] <= 16'hff01; // 0x800012cc
    mem[1204] <= 16'h0007; // 0x800012d0
    mem[1205] <= 16'h0081; // 0x800012d4
    mem[1206] <= 16'h0005; // 0x800012d8
    mem[1207] <= 16'h0011; // 0x800012dc
    mem[1208] <= 16'h0091; // 0x800012e0
    mem[1209] <= 16'h00d4; // 0x800012e4
    mem[1210] <= 16'h0047; // 0x800012e8
    mem[1211] <= 16'h0005; // 0x800012ec
    mem[1212] <= 16'h0050; // 0x800012f0
    mem[1213] <= 16'h00d4; // 0x800012f4
    mem[1214] <= 16'h0087; // 0x800012f8
    mem[1215] <= 16'h0004; // 0x800012fc
    mem[1216] <= 16'h00d4; // 0x80001300
    mem[1217] <= 16'h00c7; // 0x80001304
    mem[1218] <= 16'h00d4; // 0x80001308
    mem[1219] <= 16'h0107; // 0x8000130c
    mem[1220] <= 16'h00d4; // 0x80001310
    mem[1221] <= 16'h0147; // 0x80001314
    mem[1222] <= 16'h00d4; // 0x80001318
    mem[1223] <= 16'h0187; // 0x8000131c
    mem[1224] <= 16'h00d4; // 0x80001320
    mem[1225] <= 16'h01c7; // 0x80001324
    mem[1226] <= 16'h00d4; // 0x80001328
    mem[1227] <= 16'h0207; // 0x8000132c
    mem[1228] <= 16'h02d4; // 0x80001330
    mem[1229] <= 16'h0247; // 0x80001334
    mem[1230] <= 16'h02d4; // 0x80001338
    mem[1231] <= 16'h0287; // 0x8000133c
    mem[1232] <= 16'h02d4; // 0x80001340
    mem[1233] <= 16'h02c7; // 0x80001344
    mem[1234] <= 16'h02f4; // 0x80001348
    mem[1235] <= 16'h00e4; // 0x8000134c
    mem[1236] <= 16'h00e4; // 0x80001350
    mem[1237] <= 16'h0004; // 0x80001354
    mem[1238] <= 16'h00f4; // 0x80001358
    mem[1239] <= 16'hf39f; // 0x8000135c
    mem[1240] <= 16'h0044; // 0x80001360
    mem[1241] <= 16'h0607; // 0x80001364
    mem[1242] <= 16'h0004; // 0x80001368
    mem[1243] <= 16'h00c1; // 0x8000136c
    mem[1244] <= 16'h0081; // 0x80001370
    mem[1245] <= 16'h0007; // 0x80001374
    mem[1246] <= 16'h00e4; // 0x80001378
    mem[1247] <= 16'h0047; // 0x8000137c
    mem[1248] <= 16'h00e4; // 0x80001380
    mem[1249] <= 16'h0087; // 0x80001384
    mem[1250] <= 16'h00e4; // 0x80001388
    mem[1251] <= 16'h00c7; // 0x8000138c
    mem[1252] <= 16'h00e4; // 0x80001390
    mem[1253] <= 16'h0107; // 0x80001394
    mem[1254] <= 16'h00e4; // 0x80001398
    mem[1255] <= 16'h0147; // 0x8000139c
    mem[1256] <= 16'h00e4; // 0x800013a0
    mem[1257] <= 16'h0187; // 0x800013a4
    mem[1258] <= 16'h00e4; // 0x800013a8
    mem[1259] <= 16'h01c7; // 0x800013ac
    mem[1260] <= 16'h00e4; // 0x800013b0
    mem[1261] <= 16'h0207; // 0x800013b4
    mem[1262] <= 16'h02e4; // 0x800013b8
    mem[1263] <= 16'h0247; // 0x800013bc
    mem[1264] <= 16'h02e4; // 0x800013c0
    mem[1265] <= 16'h0287; // 0x800013c4
    mem[1266] <= 16'h02e4; // 0x800013c8
    mem[1267] <= 16'h02c7; // 0x800013cc
    mem[1268] <= 16'h02f4; // 0x800013d0
    mem[1269] <= 16'h0041; // 0x800013d4
    mem[1270] <= 16'h0101; // 0x800013d8
    mem[1271] <= 16'h0000; // 0x800013dc
    mem[1272] <= 16'h0060; // 0x800013e0
    mem[1273] <= 16'h00f4; // 0x800013e4
    mem[1274] <= 16'h0084; // 0x800013e8
    mem[1275] <= 16'h0084; // 0x800013ec
    mem[1276] <= 16'hdb1f; // 0x800013f0
    mem[1277] <= 16'h0000; // 0x800013f4
    mem[1278] <= 16'h1007; // 0x800013f8
    mem[1279] <= 16'h0007; // 0x800013fc
    mem[1280] <= 16'h00c4; // 0x80001400
    mem[1281] <= 16'h00c4; // 0x80001404
    mem[1282] <= 16'h00f4; // 0x80001408
    mem[1283] <= 16'h00c1; // 0x8000140c
    mem[1284] <= 16'h0081; // 0x80001410
    mem[1285] <= 16'h0041; // 0x80001414
    mem[1286] <= 16'h00a0; // 0x80001418
    mem[1287] <= 16'h0101; // 0x8000141c
    mem[1288] <= 16'hc29f; // 0x80001420
    mem[1289] <= 16'h0000; // 0x80001424
    mem[1290] <= 16'h0c47; // 0x80001428
    mem[1291] <= 16'h0007; // 0x8000142c
    mem[1292] <= 16'h0000; // 0x80001430
    mem[1293] <= 16'h0b57; // 0x80001434
    mem[1294] <= 16'hfbf7; // 0x80001438
    mem[1295] <= 16'h0017; // 0x8000143c
    mem[1296] <= 16'h00d7; // 0x80001440
    mem[1297] <= 16'h00f7; // 0x80001444
    mem[1298] <= 16'h0420; // 0x80001448
    mem[1299] <= 16'h0000; // 0x8000144c
    mem[1300] <= 16'h08f2; // 0x80001450
    mem[1301] <= 16'h0000; // 0x80001454
    mem[1302] <= 16'h0410; // 0x80001458
    mem[1303] <= 16'h0000; // 0x8000145c
    mem[1304] <= 16'h08f2; // 0x80001460
    mem[1305] <= 16'h0000; // 0x80001464
    mem[1306] <= 16'h0802; // 0x80001468
    mem[1307] <= 16'h0000; // 0x8000146c
    mem[1308] <= 16'h8000; // 0x80001470
    mem[1309] <= 16'h0007; // 0x80001474
    mem[1310] <= 16'hfe07; // 0x80001478
    mem[1311] <= 16'h0ff5; // 0x8000147c
    mem[1312] <= 16'h00a7; // 0x80001480
    mem[1313] <= 16'h8000; // 0x80001484
    mem[1314] <= 16'h0007; // 0x80001488
    mem[1315] <= 16'hfe07; // 0x8000148c
    mem[1316] <= 16'h0000; // 0x80001490
    mem[1317] <= 16'h0000; // 0x80001494
    mem[1318] <= 16'h0010; // 0x80001498
    mem[1319] <= 16'h0005; // 0x8000149c
    mem[1320] <= 16'h02b7; // 0x800014a0
    mem[1321] <= 16'h0005; // 0x800014a4
    mem[1322] <= 16'h0005; // 0x800014a8
    mem[1323] <= 16'h0007; // 0x800014ac
    mem[1324] <= 16'h0047; // 0x800014b0
    mem[1325] <= 16'h0000; // 0x800014b4
    mem[1326] <= 16'h00f7; // 0x800014b8
    mem[1327] <= 16'h0000; // 0x800014bc
    mem[1328] <= 16'h0047; // 0x800014c0
    mem[1329] <= 16'h00d5; // 0x800014c4
    mem[1330] <= 16'h0000; // 0x800014c8
    mem[1331] <= 16'h0007; // 0x800014cc
    mem[1332] <= 16'h0000; // 0x800014d0
    mem[1333] <= 16'h0005; // 0x800014d4
    mem[1334] <= 16'h0077; // 0x800014d8
    mem[1335] <= 16'hff87; // 0x800014dc
    mem[1336] <= 16'h0087; // 0x800014e0
    mem[1337] <= 16'h00d5; // 0x800014e4
    mem[1338] <= 16'h0047; // 0x800014e8
    mem[1339] <= 16'h0007; // 0x800014ec
    mem[1340] <= 16'h0000; // 0x800014f0
    mem[1341] <= 16'h0010; // 0x800014f4
    mem[1342] <= 16'h0005; // 0x800014f8
    mem[1343] <= 16'h00b7; // 0x800014fc
    mem[1344] <= 16'h0005; // 0x80001500
    mem[1345] <= 16'h0007; // 0x80001504
    mem[1346] <= 16'h0047; // 0x80001508
    mem[1347] <= 16'h00f7; // 0x8000150c
    mem[1348] <= 16'h41f5; // 0x80001510
    mem[1349] <= 16'h0000; // 0x80001514
    mem[1350] <= 16'h0005; // 0x80001518
    mem[1351] <= 16'h0077; // 0x8000151c
    mem[1352] <= 16'hff87; // 0x80001520
    mem[1353] <= 16'h0087; // 0x80001524
    mem[1354] <= 16'h00d5; // 0x80001528
    mem[1355] <= 16'h0047; // 0x8000152c
    mem[1356] <= 16'h0007; // 0x80001530
    mem[1357] <= 16'h0000; // 0x80001534
    mem[1358] <= 16'h0005; // 0x80001538
    mem[1359] <= 16'h00a7; // 0x8000153c
    mem[1360] <= 16'h0005; // 0x80001540
    mem[1361] <= 16'h0017; // 0x80001544
    mem[1362] <= 16'h00f5; // 0x80001548
    mem[1363] <= 16'h0000; // 0x8000154c
    mem[1364] <= 16'hed01; // 0x80001550
    mem[1365] <= 16'h1181; // 0x80001554
    mem[1366] <= 16'h0006; // 0x80001558
    mem[1367] <= 16'h0000; // 0x8000155c
    mem[1368] <= 16'h1281; // 0x80001560
    mem[1369] <= 16'h1321; // 0x80001564
    mem[1370] <= 16'h1151; // 0x80001568
    mem[1371] <= 16'h1161; // 0x8000156c
    mem[1372] <= 16'h1171; // 0x80001570
    mem[1373] <= 16'h1211; // 0x80001574
    mem[1374] <= 16'h1291; // 0x80001578
    mem[1375] <= 16'h1131; // 0x8000157c
    mem[1376] <= 16'h1141; // 0x80001580
    mem[1377] <= 16'h0005; // 0x80001584
    mem[1378] <= 16'h0005; // 0x80001588
    mem[1379] <= 16'h0006; // 0x8000158c
    mem[1380] <= 16'h0007; // 0x80001590
    mem[1381] <= 16'h6640; // 0x80001594
    mem[1382] <= 16'h00a1; // 0x80001598
    mem[1383] <= 16'h0000; // 0x8000159c
    mem[1384] <= 16'h0e04; // 0x800015a0
    mem[1385] <= 16'h0041; // 0x800015a4
    mem[1386] <= 16'h0010; // 0x800015a8
    mem[1387] <= 16'h000a; // 0x800015ac
    mem[1388] <= 16'h0000; // 0x800015b0
    mem[1389] <= 16'h0009; // 0x800015b4
    mem[1390] <= 16'h0004; // 0x800015b8
    mem[1391] <= 16'h1c80; // 0x800015bc
    mem[1392] <= 16'h000a; // 0x800015c0
    mem[1393] <= 16'h0000; // 0x800015c4
    mem[1394] <= 16'h0005; // 0x800015c8
    mem[1395] <= 16'h0005; // 0x800015cc
    mem[1396] <= 16'h6280; // 0x800015d0
    mem[1397] <= 16'h00a9; // 0x800015d4
    mem[1398] <= 16'h0014; // 0x800015d8
    mem[1399] <= 16'h0049; // 0x800015dc
    mem[1400] <= 16'h008b; // 0x800015e0
    mem[1401] <= 16'h000a; // 0x800015e4
    mem[1402] <= 16'hfc5f; // 0x800015e8
    mem[1403] <= 16'hff59; // 0x800015ec
    mem[1404] <= 16'hfffc; // 0x800015f0
    mem[1405] <= 16'h038a; // 0x800015f4
    mem[1406] <= 16'h0000; // 0x800015f8
    mem[1407] <= 16'h000b; // 0x800015fc
    mem[1408] <= 16'hfff4; // 0x80001600
    mem[1409] <= 16'he6df; // 0x80001604
    mem[1410] <= 16'h0014; // 0x80001608
    mem[1411] <= 16'hfefa; // 0x8000160c
    mem[1412] <= 16'h0540; // 0x80001610
    mem[1413] <= 16'h0024; // 0x80001614
    mem[1414] <= 16'h0081; // 0x80001618
    mem[1415] <= 16'h0090; // 0x8000161c
    mem[1416] <= 16'h0300; // 0x80001620
    mem[1417] <= 16'h0570; // 0x80001624
    mem[1418] <= 16'h0004; // 0x80001628
    mem[1419] <= 16'h0000; // 0x8000162c
    mem[1420] <= 16'hfff4; // 0x80001630
    mem[1421] <= 16'h0009; // 0x80001634
    mem[1422] <= 16'h00f9; // 0x80001638
    mem[1423] <= 16'h000a; // 0x8000163c
    mem[1424] <= 16'h00a7; // 0x80001640
    mem[1425] <= 16'he2df; // 0x80001644
    mem[1426] <= 16'h0014; // 0x80001648
    mem[1427] <= 16'hffc4; // 0x8000164c
    mem[1428] <= 16'hfcf0; // 0x80001650
    mem[1429] <= 16'h12c1; // 0x80001654
    mem[1430] <= 16'h1281; // 0x80001658
    mem[1431] <= 16'h1241; // 0x8000165c
    mem[1432] <= 16'h1201; // 0x80001660
    mem[1433] <= 16'h11c1; // 0x80001664
    mem[1434] <= 16'h1181; // 0x80001668
    mem[1435] <= 16'h1141; // 0x8000166c
    mem[1436] <= 16'h1101; // 0x80001670
    mem[1437] <= 16'h10c1; // 0x80001674
    mem[1438] <= 16'h1081; // 0x80001678
    mem[1439] <= 16'h1301; // 0x8000167c
    mem[1440] <= 16'h0000; // 0x80001680
    mem[1441] <= 16'hf359; // 0x80001684
    mem[1442] <= 16'h0010; // 0x80001688
    mem[1443] <= 16'hfffc; // 0x8000168c
    mem[1444] <= 16'h0000; // 0x80001690
    mem[1445] <= 16'hf78a; // 0x80001694
    mem[1446] <= 16'hf7df; // 0x80001698
    mem[1447] <= 16'hed01; // 0x8000169c
    mem[1448] <= 16'h1281; // 0x800016a0
    mem[1449] <= 16'h1321; // 0x800016a4
    mem[1450] <= 16'h0006; // 0x800016a8
    mem[1451] <= 16'h0006; // 0x800016ac
    mem[1452] <= 16'h1141; // 0x800016b0
    mem[1453] <= 16'h0007; // 0x800016b4
    mem[1454] <= 16'h0005; // 0x800016b8
    mem[1455] <= 16'h0000; // 0x800016bc
    mem[1456] <= 16'h0009; // 0x800016c0
    mem[1457] <= 16'h0004; // 0x800016c4
    mem[1458] <= 16'h1161; // 0x800016c8
    mem[1459] <= 16'h1171; // 0x800016cc
    mem[1460] <= 16'h1181; // 0x800016d0
    mem[1461] <= 16'h1191; // 0x800016d4
    mem[1462] <= 16'h1211; // 0x800016d8
    mem[1463] <= 16'h1291; // 0x800016dc
    mem[1464] <= 16'h1131; // 0x800016e0
    mem[1465] <= 16'h1151; // 0x800016e4
    mem[1466] <= 16'h0007; // 0x800016e8
    mem[1467] <= 16'h0007; // 0x800016ec
    mem[1468] <= 16'h0008; // 0x800016f0
    mem[1469] <= 16'h5040; // 0x800016f4
    mem[1470] <= 16'h00a1; // 0x800016f8
    mem[1471] <= 16'h0000; // 0x800016fc
    mem[1472] <= 16'h0e04; // 0x80001700
    mem[1473] <= 16'h0041; // 0x80001704
    mem[1474] <= 16'h0010; // 0x80001708
    mem[1475] <= 16'h000b; // 0x8000170c
    mem[1476] <= 16'h0000; // 0x80001710
    mem[1477] <= 16'h0009; // 0x80001714
    mem[1478] <= 16'h0004; // 0x80001718
    mem[1479] <= 16'h0680; // 0x8000171c
    mem[1480] <= 16'h000b; // 0x80001720
    mem[1481] <= 16'h0000; // 0x80001724
    mem[1482] <= 16'h0005; // 0x80001728
    mem[1483] <= 16'h0005; // 0x8000172c
    mem[1484] <= 16'h4c80; // 0x80001730
    mem[1485] <= 16'h00a9; // 0x80001734
    mem[1486] <= 16'h0014; // 0x80001738
    mem[1487] <= 16'h0049; // 0x8000173c
    mem[1488] <= 16'h008b; // 0x80001740
    mem[1489] <= 16'h000a; // 0x80001744
    mem[1490] <= 16'hfc5f; // 0x80001748
    mem[1491] <= 16'hff69; // 0x8000174c
    mem[1492] <= 16'hfffc; // 0x80001750
    mem[1493] <= 16'h039a; // 0x80001754
    mem[1494] <= 16'h000a; // 0x80001758
    mem[1495] <= 16'h000c; // 0x8000175c
    mem[1496] <= 16'hfff4; // 0x80001760
    mem[1497] <= 16'hdd5f; // 0x80001764
    mem[1498] <= 16'h0014; // 0x80001768
    mem[1499] <= 16'hfefa; // 0x8000176c
    mem[1500] <= 16'h0550; // 0x80001770
    mem[1501] <= 16'h0024; // 0x80001774
    mem[1502] <= 16'h0081; // 0x80001778
    mem[1503] <= 16'h0090; // 0x8000177c
    mem[1504] <= 16'h0300; // 0x80001780
    mem[1505] <= 16'h0570; // 0x80001784
    mem[1506] <= 16'h0004; // 0x80001788
    mem[1507] <= 16'h000a; // 0x8000178c
    mem[1508] <= 16'hfff4; // 0x80001790
    mem[1509] <= 16'h0009; // 0x80001794
    mem[1510] <= 16'h00f9; // 0x80001798
    mem[1511] <= 16'h000a; // 0x8000179c
    mem[1512] <= 16'h00a7; // 0x800017a0
    mem[1513] <= 16'hd95f; // 0x800017a4
    mem[1514] <= 16'h0014; // 0x800017a8
    mem[1515] <= 16'hffc4; // 0x800017ac
    mem[1516] <= 16'hfcf0; // 0x800017b0
    mem[1517] <= 16'h12c1; // 0x800017b4
    mem[1518] <= 16'h1281; // 0x800017b8
    mem[1519] <= 16'h1241; // 0x800017bc
    mem[1520] <= 16'h1201; // 0x800017c0
    mem[1521] <= 16'h11c1; // 0x800017c4
    mem[1522] <= 16'h1181; // 0x800017c8
    mem[1523] <= 16'h1141; // 0x800017cc
    mem[1524] <= 16'h1101; // 0x800017d0
    mem[1525] <= 16'h10c1; // 0x800017d4
    mem[1526] <= 16'h1081; // 0x800017d8
    mem[1527] <= 16'h1041; // 0x800017dc
    mem[1528] <= 16'h1301; // 0x800017e0
    mem[1529] <= 16'h0000; // 0x800017e4
    mem[1530] <= 16'hf169; // 0x800017e8
    mem[1531] <= 16'h0010; // 0x800017ec
    mem[1532] <= 16'hfffc; // 0x800017f0
    mem[1533] <= 16'h0000; // 0x800017f4
    mem[1534] <= 16'hf79a; // 0x800017f8
    mem[1535] <= 16'hf79f; // 0x800017fc
    mem[1536] <= 16'hb000; // 0x80001800
    mem[1537] <= 16'h0205; // 0x80001804
    mem[1538] <= 16'h0000; // 0x80001808
    mem[1539] <= 16'hcf87; // 0x8000180c
    mem[1540] <= 16'h40e7; // 0x80001810
    mem[1541] <= 16'h0000; // 0x80001814
    mem[1542] <= 16'hc2c7; // 0x80001818
    mem[1543] <= 16'h0000; // 0x8000181c
    mem[1544] <= 16'hcce2; // 0x80001820
    mem[1545] <= 16'h0000; // 0x80001824
    mem[1546] <= 16'hcdc7; // 0x80001828
    mem[1547] <= 16'h00f7; // 0x8000182c
    mem[1548] <= 16'hb020; // 0x80001830
    mem[1549] <= 16'h0205; // 0x80001834
    mem[1550] <= 16'h0000; // 0x80001838
    mem[1551] <= 16'hccc6; // 0x8000183c
    mem[1552] <= 16'h40d7; // 0x80001840
    mem[1553] <= 16'h0000; // 0x80001844
    mem[1554] <= 16'hc046; // 0x80001848
    mem[1555] <= 16'h0000; // 0x8000184c
    mem[1556] <= 16'hcad2; // 0x80001850
    mem[1557] <= 16'h00f7; // 0x80001854
    mem[1558] <= 16'h0000; // 0x80001858
    mem[1559] <= 16'h0015; // 0x8000185c
    mem[1560] <= 16'hffff; // 0x80001860
    mem[1561] <= 16'h7a06; // 0x80001864
    mem[1562] <= 16'h0015; // 0x80001868
    mem[1563] <= 16'h0000; // 0x8000186c
    mem[1564] <= 16'h00e6; // 0x80001870
    mem[1565] <= 16'h00f6; // 0x80001874
    mem[1566] <= 16'h0000; // 0x80001878
    mem[1567] <= 16'hff01; // 0x8000187c
    mem[1568] <= 16'h5390; // 0x80001880
    mem[1569] <= 16'h0011; // 0x80001884
    mem[1570] <= 16'hfd5f; // 0x80001888
    mem[1571] <= 16'hff01; // 0x8000188c
    mem[1572] <= 16'h0011; // 0x80001890
    mem[1573] <= 16'hfc9f; // 0x80001894
    mem[1574] <= 16'hff01; // 0x80001898
    mem[1575] <= 16'h0860; // 0x8000189c
    mem[1576] <= 16'h0011; // 0x800018a0
    mem[1577] <= 16'hfe9f; // 0x800018a4
    mem[1578] <= 16'h0005; // 0x800018a8
    mem[1579] <= 16'h0000; // 0x800018ac
    mem[1580] <= 16'h0000; // 0x800018b0
    mem[1581] <= 16'h00c5; // 0x800018b4
    mem[1582] <= 16'h00a7; // 0x800018b8
    mem[1583] <= 16'h0037; // 0x800018bc
    mem[1584] <= 16'h0a07; // 0x800018c0
    mem[1585] <= 16'h00c5; // 0x800018c4
    mem[1586] <= 16'h0f05; // 0x800018c8
    mem[1587] <= 16'h0045; // 0x800018cc
    mem[1588] <= 16'h0045; // 0x800018d0
    mem[1589] <= 16'h00e5; // 0x800018d4
    mem[1590] <= 16'h00d5; // 0x800018d8
    mem[1591] <= 16'h00b5; // 0x800018dc
    mem[1592] <= 16'h0017; // 0x800018e0
    mem[1593] <= 16'h0016; // 0x800018e4
    mem[1594] <= 16'h0037; // 0x800018e8
    mem[1595] <= 16'h00d7; // 0x800018ec
    mem[1596] <= 16'h0017; // 0x800018f0
    mem[1597] <= 16'h00e7; // 0x800018f4
    mem[1598] <= 16'h0807; // 0x800018f8
    mem[1599] <= 16'h00a6; // 0x800018fc
    mem[1600] <= 16'h0807; // 0x80001900
    mem[1601] <= 16'hffc6; // 0x80001904
    mem[1602] <= 16'h0027; // 0x80001908
    mem[1603] <= 16'h0017; // 0x8000190c
    mem[1604] <= 16'h0027; // 0x80001910
    mem[1605] <= 16'h0005; // 0x80001914
    mem[1606] <= 16'h0005; // 0x80001918
    mem[1607] <= 16'h0000; // 0x8000191c
    mem[1608] <= 16'h0006; // 0x80001920
    mem[1609] <= 16'h0017; // 0x80001924
    mem[1610] <= 16'h0046; // 0x80001928
    mem[1611] <= 16'h01c8; // 0x8000192c
    mem[1612] <= 16'h0048; // 0x80001930
    mem[1613] <= 16'hfef7; // 0x80001934
    mem[1614] <= 16'h0065; // 0x80001938
    mem[1615] <= 16'h0065; // 0x8000193c
    mem[1616] <= 16'h0666; // 0x80001940
    mem[1617] <= 16'h0005; // 0x80001944
    mem[1618] <= 16'h0017; // 0x80001948
    mem[1619] <= 16'h00d7; // 0x8000194c
    mem[1620] <= 16'h0507; // 0x80001950
    mem[1621] <= 16'h0015; // 0x80001954
    mem[1622] <= 16'h0027; // 0x80001958
    mem[1623] <= 16'h00d7; // 0x8000195c
    mem[1624] <= 16'h0507; // 0x80001960
    mem[1625] <= 16'h0025; // 0x80001964
    mem[1626] <= 16'h00e7; // 0x80001968
    mem[1627] <= 16'h0000; // 0x8000196c
    mem[1628] <= 16'h00c5; // 0x80001970
    mem[1629] <= 16'h02c5; // 0x80001974
    mem[1630] <= 16'h0005; // 0x80001978
    mem[1631] <= 16'h0045; // 0x8000197c
    mem[1632] <= 16'hffc5; // 0x80001980
    mem[1633] <= 16'h0047; // 0x80001984
    mem[1634] <= 16'hfee7; // 0x80001988
    mem[1635] <= 16'hfec7; // 0x8000198c
    mem[1636] <= 16'h0000; // 0x80001990
    mem[1637] <= 16'h0005; // 0x80001994
    mem[1638] <= 16'h0015; // 0x80001998
    mem[1639] <= 16'hfff5; // 0x8000199c
    mem[1640] <= 16'h0017; // 0x800019a0
    mem[1641] <= 16'hfee7; // 0x800019a4
    mem[1642] <= 16'hfef8; // 0x800019a8
    mem[1643] <= 16'h0000; // 0x800019ac
    mem[1644] <= 16'h0000; // 0x800019b0
    mem[1645] <= 16'h0000; // 0x800019b4
    mem[1646] <= 16'hff01; // 0x800019b8
    mem[1647] <= 16'h00c5; // 0x800019bc
    mem[1648] <= 16'h0081; // 0x800019c0
    mem[1649] <= 16'h0011; // 0x800019c4
    mem[1650] <= 16'h0037; // 0x800019c8
    mem[1651] <= 16'h0005; // 0x800019cc
    mem[1652] <= 16'h0207; // 0x800019d0
    mem[1653] <= 16'h00c5; // 0x800019d4
    mem[1654] <= 16'h00c5; // 0x800019d8
    mem[1655] <= 16'h40a6; // 0x800019dc
    mem[1656] <= 16'h0ff5; // 0x800019e0
    mem[1657] <= 16'hfd5f; // 0x800019e4
    mem[1658] <= 16'h00c1; // 0x800019e8
    mem[1659] <= 16'h0004; // 0x800019ec
    mem[1660] <= 16'h0081; // 0x800019f0
    mem[1661] <= 16'h0101; // 0x800019f4
    mem[1662] <= 16'h0000; // 0x800019f8
    mem[1663] <= 16'h0ff5; // 0x800019fc
    mem[1664] <= 16'h0087; // 0x80001a00
    mem[1665] <= 16'h00b7; // 0x80001a04
    mem[1666] <= 16'h0107; // 0x80001a08
    mem[1667] <= 16'h00c5; // 0x80001a0c
    mem[1668] <= 16'h00f7; // 0x80001a10
    mem[1669] <= 16'hfcc5; // 0x80001a14
    mem[1670] <= 16'h0005; // 0x80001a18
    mem[1671] <= 16'h0047; // 0x80001a1c
    mem[1672] <= 16'hfee7; // 0x80001a20
    mem[1673] <= 16'hfec7; // 0x80001a24
    mem[1674] <= 16'h00c1; // 0x80001a28
    mem[1675] <= 16'h0004; // 0x80001a2c
    mem[1676] <= 16'h0081; // 0x80001a30
    mem[1677] <= 16'h0101; // 0x80001a34
    mem[1678] <= 16'h0000; // 0x80001a38
    mem[1679] <= 16'hff01; // 0x80001a3c
    mem[1680] <= 16'h0081; // 0x80001a40
    mem[1681] <= 16'h0091; // 0x80001a44
    mem[1682] <= 16'h0002; // 0x80001a48
    mem[1683] <= 16'h0002; // 0x80001a4c
    mem[1684] <= 16'h4084; // 0x80001a50
    mem[1685] <= 16'h0004; // 0x80001a54
    mem[1686] <= 16'h0000; // 0x80001a58
    mem[1687] <= 16'h2885; // 0x80001a5c
    mem[1688] <= 16'h0002; // 0x80001a60
    mem[1689] <= 16'h0011; // 0x80001a64
    mem[1690] <= 16'h0121; // 0x80001a68
    mem[1691] <= 16'h0002; // 0x80001a6c
    mem[1692] <= 16'he45f; // 0x80001a70
    mem[1693] <= 16'h0002; // 0x80001a74
    mem[1694] <= 16'h0089; // 0x80001a78
    mem[1695] <= 16'h4096; // 0x80001a7c
    mem[1696] <= 16'h00c1; // 0x80001a80
    mem[1697] <= 16'h0081; // 0x80001a84
    mem[1698] <= 16'h0041; // 0x80001a88
    mem[1699] <= 16'h0001; // 0x80001a8c
    mem[1700] <= 16'h0000; // 0x80001a90
    mem[1701] <= 16'h0101; // 0x80001a94
    mem[1702] <= 16'hf21f; // 0x80001a98
    mem[1703] <= 16'h0005; // 0x80001a9c
    mem[1704] <= 16'h0007; // 0x80001aa0
    mem[1705] <= 16'h0005; // 0x80001aa4
    mem[1706] <= 16'h0017; // 0x80001aa8
    mem[1707] <= 16'h0007; // 0x80001aac
    mem[1708] <= 16'hfe07; // 0x80001ab0
    mem[1709] <= 16'h40a7; // 0x80001ab4
    mem[1710] <= 16'h0000; // 0x80001ab8
    mem[1711] <= 16'h0000; // 0x80001abc
    mem[1712] <= 16'h0000; // 0x80001ac0
    mem[1713] <= 16'hfe01; // 0x80001ac4
    mem[1714] <= 16'h0131; // 0x80001ac8
    mem[1715] <= 16'h0005; // 0x80001acc
    mem[1716] <= 16'h0121; // 0x80001ad0
    mem[1717] <= 16'h0005; // 0x80001ad4
    mem[1718] <= 16'h0009; // 0x80001ad8
    mem[1719] <= 16'h0081; // 0x80001adc
    mem[1720] <= 16'h0091; // 0x80001ae0
    mem[1721] <= 16'h0011; // 0x80001ae4
    mem[1722] <= 16'h0000; // 0x80001ae8
    mem[1723] <= 16'h8000; // 0x80001aec
    mem[1724] <= 16'hfadf; // 0x80001af0
    mem[1725] <= 16'h02a4; // 0x80001af4
    mem[1726] <= 16'h0004; // 0x80001af8
    mem[1727] <= 16'hfe07; // 0x80001afc
    mem[1728] <= 16'h0009; // 0x80001b00
    mem[1729] <= 16'h00f4; // 0x80001b04
    mem[1730] <= 16'h0004; // 0x80001b08
    mem[1731] <= 16'hfe07; // 0x80001b0c
    mem[1732] <= 16'h0009; // 0x80001b10
    mem[1733] <= 16'h0014; // 0x80001b14
    mem[1734] <= 16'h0019; // 0x80001b18
    mem[1735] <= 16'hf81f; // 0x80001b1c
    mem[1736] <= 16'hfca4; // 0x80001b20
    mem[1737] <= 16'h01c1; // 0x80001b24
    mem[1738] <= 16'h0181; // 0x80001b28
    mem[1739] <= 16'h0141; // 0x80001b2c
    mem[1740] <= 16'h0101; // 0x80001b30
    mem[1741] <= 16'h00c1; // 0x80001b34
    mem[1742] <= 16'h0201; // 0x80001b38
    mem[1743] <= 16'h0000; // 0x80001b3c
    mem[1744] <= 16'hfd01; // 0x80001b40
    mem[1745] <= 16'h0211; // 0x80001b44
    mem[1746] <= 16'h00f5; // 0x80001b48
    mem[1747] <= 16'h0090; // 0x80001b4c
    mem[1748] <= 16'h0300; // 0x80001b50
    mem[1749] <= 16'h00f6; // 0x80001b54
    mem[1750] <= 16'h0570; // 0x80001b58
    mem[1751] <= 16'h00e7; // 0x80001b5c
    mem[1752] <= 16'h0045; // 0x80001b60
    mem[1753] <= 16'h00e1; // 0x80001b64
    mem[1754] <= 16'h00f7; // 0x80001b68
    mem[1755] <= 16'h0090; // 0x80001b6c
    mem[1756] <= 16'h0570; // 0x80001b70
    mem[1757] <= 16'h00f6; // 0x80001b74
    mem[1758] <= 16'h0300; // 0x80001b78
    mem[1759] <= 16'h00e7; // 0x80001b7c
    mem[1760] <= 16'h0085; // 0x80001b80
    mem[1761] <= 16'h00e1; // 0x80001b84
    mem[1762] <= 16'h00f7; // 0x80001b88
    mem[1763] <= 16'h0090; // 0x80001b8c
    mem[1764] <= 16'h0570; // 0x80001b90
    mem[1765] <= 16'h00f6; // 0x80001b94
    mem[1766] <= 16'h0300; // 0x80001b98
    mem[1767] <= 16'h00e7; // 0x80001b9c
    mem[1768] <= 16'h00c5; // 0x80001ba0
    mem[1769] <= 16'h00e1; // 0x80001ba4
    mem[1770] <= 16'h00f7; // 0x80001ba8
    mem[1771] <= 16'h0090; // 0x80001bac
    mem[1772] <= 16'h0570; // 0x80001bb0
    mem[1773] <= 16'h00f6; // 0x80001bb4
    mem[1774] <= 16'h0300; // 0x80001bb8
    mem[1775] <= 16'h00e7; // 0x80001bbc
    mem[1776] <= 16'h0105; // 0x80001bc0
    mem[1777] <= 16'h00e1; // 0x80001bc4
    mem[1778] <= 16'h00f7; // 0x80001bc8
    mem[1779] <= 16'h0090; // 0x80001bcc
    mem[1780] <= 16'h0570; // 0x80001bd0
    mem[1781] <= 16'h00f6; // 0x80001bd4
    mem[1782] <= 16'h0300; // 0x80001bd8
    mem[1783] <= 16'h00e7; // 0x80001bdc
    mem[1784] <= 16'h0145; // 0x80001be0
    mem[1785] <= 16'h00e1; // 0x80001be4
    mem[1786] <= 16'h00f7; // 0x80001be8
    mem[1787] <= 16'h0090; // 0x80001bec
    mem[1788] <= 16'h0570; // 0x80001bf0
    mem[1789] <= 16'h00f6; // 0x80001bf4
    mem[1790] <= 16'h0300; // 0x80001bf8
    mem[1791] <= 16'h00e7; // 0x80001bfc
    mem[1792] <= 16'h0185; // 0x80001c00
    mem[1793] <= 16'h00e1; // 0x80001c04
    mem[1794] <= 16'h00f7; // 0x80001c08
    mem[1795] <= 16'h0090; // 0x80001c0c
    mem[1796] <= 16'h0570; // 0x80001c10
    mem[1797] <= 16'h00f6; // 0x80001c14
    mem[1798] <= 16'h0300; // 0x80001c18
    mem[1799] <= 16'h00e7; // 0x80001c1c
    mem[1800] <= 16'h00f1; // 0x80001c20
    mem[1801] <= 16'h01c5; // 0x80001c24
    mem[1802] <= 16'h0090; // 0x80001c28
    mem[1803] <= 16'h0570; // 0x80001c2c
    mem[1804] <= 16'h00a7; // 0x80001c30
    mem[1805] <= 16'h0300; // 0x80001c34
    mem[1806] <= 16'h00f5; // 0x80001c38
    mem[1807] <= 16'h00a1; // 0x80001c3c
    mem[1808] <= 16'h00f5; // 0x80001c40
    mem[1809] <= 16'h0090; // 0x80001c44
    mem[1810] <= 16'h0570; // 0x80001c48
    mem[1811] <= 16'h00f6; // 0x80001c4c
    mem[1812] <= 16'h0300; // 0x80001c50
    mem[1813] <= 16'h00e7; // 0x80001c54
    mem[1814] <= 16'h0045; // 0x80001c58
    mem[1815] <= 16'h00e1; // 0x80001c5c
    mem[1816] <= 16'h00f7; // 0x80001c60
    mem[1817] <= 16'h0090; // 0x80001c64
    mem[1818] <= 16'h0570; // 0x80001c68
    mem[1819] <= 16'h00f6; // 0x80001c6c
    mem[1820] <= 16'h0300; // 0x80001c70
    mem[1821] <= 16'h00e7; // 0x80001c74
    mem[1822] <= 16'h0085; // 0x80001c78
    mem[1823] <= 16'h00e1; // 0x80001c7c
    mem[1824] <= 16'h00f7; // 0x80001c80
    mem[1825] <= 16'h0090; // 0x80001c84
    mem[1826] <= 16'h0570; // 0x80001c88
    mem[1827] <= 16'h00f6; // 0x80001c8c
    mem[1828] <= 16'h0300; // 0x80001c90
    mem[1829] <= 16'h00e7; // 0x80001c94
    mem[1830] <= 16'h00c5; // 0x80001c98
    mem[1831] <= 16'h00e1; // 0x80001c9c
    mem[1832] <= 16'h00f7; // 0x80001ca0
    mem[1833] <= 16'h0090; // 0x80001ca4
    mem[1834] <= 16'h0570; // 0x80001ca8
    mem[1835] <= 16'h00f6; // 0x80001cac
    mem[1836] <= 16'h0300; // 0x80001cb0
    mem[1837] <= 16'h00e7; // 0x80001cb4
    mem[1838] <= 16'h0105; // 0x80001cb8
    mem[1839] <= 16'h00e1; // 0x80001cbc
    mem[1840] <= 16'h00f7; // 0x80001cc0
    mem[1841] <= 16'h0090; // 0x80001cc4
    mem[1842] <= 16'h0570; // 0x80001cc8
    mem[1843] <= 16'h00f6; // 0x80001ccc
    mem[1844] <= 16'h0300; // 0x80001cd0
    mem[1845] <= 16'h00e7; // 0x80001cd4
    mem[1846] <= 16'h0145; // 0x80001cd8
    mem[1847] <= 16'h00e1; // 0x80001cdc
    mem[1848] <= 16'h00f7; // 0x80001ce0
    mem[1849] <= 16'h0090; // 0x80001ce4
    mem[1850] <= 16'h0570; // 0x80001ce8
    mem[1851] <= 16'h00f6; // 0x80001cec
    mem[1852] <= 16'h0300; // 0x80001cf0
    mem[1853] <= 16'h00e7; // 0x80001cf4
    mem[1854] <= 16'h0185; // 0x80001cf8
    mem[1855] <= 16'h00e1; // 0x80001cfc
    mem[1856] <= 16'h00f7; // 0x80001d00
    mem[1857] <= 16'h0090; // 0x80001d04
    mem[1858] <= 16'h0570; // 0x80001d08
    mem[1859] <= 16'h00f6; // 0x80001d0c
    mem[1860] <= 16'h0300; // 0x80001d10
    mem[1861] <= 16'h00e7; // 0x80001d14
    mem[1862] <= 16'h00f1; // 0x80001d18
    mem[1863] <= 16'h01c5; // 0x80001d1c
    mem[1864] <= 16'h0090; // 0x80001d20
    mem[1865] <= 16'h0570; // 0x80001d24
    mem[1866] <= 16'h00b7; // 0x80001d28
    mem[1867] <= 16'h0300; // 0x80001d2c
    mem[1868] <= 16'h00f5; // 0x80001d30
    mem[1869] <= 16'h00c1; // 0x80001d34
    mem[1870] <= 16'h00b1; // 0x80001d38
    mem[1871] <= 16'h0001; // 0x80001d3c
    mem[1872] <= 16'hd85f; // 0x80001d40
    mem[1873] <= 16'h02c1; // 0x80001d44
    mem[1874] <= 16'h0301; // 0x80001d48
    mem[1875] <= 16'h0000; // 0x80001d4c
    mem[1876] <= 16'h0205; // 0x80001d50
    mem[1877] <= 16'h0005; // 0x80001d54
    mem[1878] <= 16'h0207; // 0x80001d58
    mem[1879] <= 16'h00b5; // 0x80001d5c
    mem[1880] <= 16'h0005; // 0x80001d60
    mem[1881] <= 16'h00c0; // 0x80001d64
    mem[1882] <= 16'h0007; // 0x80001d68
    mem[1883] <= 16'h0007; // 0x80001d6c
    mem[1884] <= 16'h0017; // 0x80001d70
    mem[1885] <= 16'hfeb7; // 0x80001d74
    mem[1886] <= 16'h40a7; // 0x80001d78
    mem[1887] <= 16'h0000; // 0x80001d7c
    mem[1888] <= 16'h0000; // 0x80001d80
    mem[1889] <= 16'h0000; // 0x80001d84
    mem[1890] <= 16'hfc01; // 0x80001d88
    mem[1891] <= 16'h0281; // 0x80001d8c
    mem[1892] <= 16'h0321; // 0x80001d90
    mem[1893] <= 16'h0331; // 0x80001d94
    mem[1894] <= 16'h0341; // 0x80001d98
    mem[1895] <= 16'h0351; // 0x80001d9c
    mem[1896] <= 16'h0361; // 0x80001da0
    mem[1897] <= 16'h0211; // 0x80001da4
    mem[1898] <= 16'h0291; // 0x80001da8
    mem[1899] <= 16'h0171; // 0x80001dac
    mem[1900] <= 16'h0181; // 0x80001db0
    mem[1901] <= 16'h0191; // 0x80001db4
    mem[1902] <= 16'h01a1; // 0x80001db8
    mem[1903] <= 16'h0005; // 0x80001dbc
    mem[1904] <= 16'h0005; // 0x80001dc0
    mem[1905] <= 16'h00c1; // 0x80001dc4
    mem[1906] <= 16'h0000; // 0x80001dc8
    mem[1907] <= 16'h2c89; // 0x80001dcc
    mem[1908] <= 16'h0010; // 0x80001dd0
    mem[1909] <= 16'h0300; // 0x80001dd4
    mem[1910] <= 16'hfff0; // 0x80001dd8
    mem[1911] <= 16'h0004; // 0x80001ddc
    mem[1912] <= 16'h0250; // 0x80001de0
    mem[1913] <= 16'h0095; // 0x80001de4
    mem[1914] <= 16'h0605; // 0x80001de8
    mem[1915] <= 16'h0009; // 0x80001dec
    mem[1916] <= 16'h0014; // 0x80001df0
    mem[1917] <= 16'hf44f; // 0x80001df4
    mem[1918] <= 16'h0004; // 0x80001df8
    mem[1919] <= 16'hfe95; // 0x80001dfc
    mem[1920] <= 16'h00c1; // 0x80001e00
    mem[1921] <= 16'h0014; // 0x80001e04
    mem[1922] <= 16'h0014; // 0x80001e08
    mem[1923] <= 16'hfff0; // 0x80001e0c
    mem[1924] <= 16'h0006; // 0x80001e10
    mem[1925] <= 16'h000c; // 0x80001e14
    mem[1926] <= 16'h0000; // 0x80001e18
    mem[1927] <= 16'h0200; // 0x80001e1c
    mem[1928] <= 16'h0004; // 0x80001e20
    mem[1929] <= 16'h0000; // 0x80001e24
    mem[1930] <= 16'h0550; // 0x80001e28
    mem[1931] <= 16'h0090; // 0x80001e2c
    mem[1932] <= 16'h02d0; // 0x80001e30
    mem[1933] <= 16'hfdde; // 0x80001e34
    mem[1934] <= 16'h0ff7; // 0x80001e38
    mem[1935] <= 16'h0017; // 0x80001e3c
    mem[1936] <= 16'h28e6; // 0x80001e40
    mem[1937] <= 16'h0027; // 0x80001e44
    mem[1938] <= 16'h0137; // 0x80001e48
    mem[1939] <= 16'h0007; // 0x80001e4c
    mem[1940] <= 16'h0137; // 0x80001e50
    mem[1941] <= 16'h0007; // 0x80001e54
    mem[1942] <= 16'h03c1; // 0x80001e58
    mem[1943] <= 16'h0381; // 0x80001e5c
    mem[1944] <= 16'h0341; // 0x80001e60
    mem[1945] <= 16'h0301; // 0x80001e64
    mem[1946] <= 16'h02c1; // 0x80001e68
    mem[1947] <= 16'h0281; // 0x80001e6c
    mem[1948] <= 16'h0241; // 0x80001e70
    mem[1949] <= 16'h0201; // 0x80001e74
    mem[1950] <= 16'h01c1; // 0x80001e78
    mem[1951] <= 16'h0181; // 0x80001e7c
    mem[1952] <= 16'h0141; // 0x80001e80
    mem[1953] <= 16'h0101; // 0x80001e84
    mem[1954] <= 16'h0401; // 0x80001e88
    mem[1955] <= 16'h0000; // 0x80001e8c
    mem[1956] <= 16'h000c; // 0x80001e90
    mem[1957] <= 16'h0000; // 0x80001e94
    mem[1958] <= 16'h0017; // 0x80001e98
    mem[1959] <= 16'h0004; // 0x80001e9c
    mem[1960] <= 16'hf95f; // 0x80001ea0
    mem[1961] <= 16'h2a08; // 0x80001ea4
    mem[1962] <= 16'h0100; // 0x80001ea8
    mem[1963] <= 16'h00c1; // 0x80001eac
    mem[1964] <= 16'hde8f; // 0x80001eb0
    mem[1965] <= 16'h0005; // 0x80001eb4
    mem[1966] <= 16'h0005; // 0x80001eb8
    mem[1967] <= 16'h000b; // 0x80001ebc
    mem[1968] <= 16'h000c; // 0x80001ec0
    mem[1969] <= 16'h0004; // 0x80001ec4
    mem[1970] <= 16'h0009; // 0x80001ec8
    mem[1971] <= 16'hfd0f; // 0x80001ecc
    mem[1972] <= 16'hf0df; // 0x80001ed0
    mem[1973] <= 16'h2808; // 0x80001ed4
    mem[1974] <= 16'h0009; // 0x80001ed8
    mem[1975] <= 16'h0250; // 0x80001edc
    mem[1976] <= 16'he58f; // 0x80001ee0
    mem[1977] <= 16'hef9f; // 0x80001ee4
    mem[1978] <= 16'h0008; // 0x80001ee8
    mem[1979] <= 16'h0017; // 0x80001eec
    mem[1980] <= 16'h0048; // 0x80001ef0
    mem[1981] <= 16'h0004; // 0x80001ef4
    mem[1982] <= 16'h000b; // 0x80001ef8
    mem[1983] <= 16'hf20c; // 0x80001efc
    mem[1984] <= 16'h0004; // 0x80001f00
    mem[1985] <= 16'hfff0; // 0x80001f04
    mem[1986] <= 16'hf2df; // 0x80001f08
    mem[1987] <= 16'h0017; // 0x80001f0c
    mem[1988] <= 16'h0003; // 0x80001f10
    mem[1989] <= 16'h0004; // 0x80001f14
    mem[1990] <= 16'hf1df; // 0x80001f18
    mem[1991] <= 16'h0017; // 0x80001f1c
    mem[1992] <= 16'h000a; // 0x80001f20
    mem[1993] <= 16'h0004; // 0x80001f24
    mem[1994] <= 16'hf0df; // 0x80001f28
    mem[1995] <= 16'h0017; // 0x80001f2c
    mem[1996] <= 16'hfd0e; // 0x80001f30
    mem[1997] <= 16'hfd0e; // 0x80001f34
    mem[1998] <= 16'h1cf5; // 0x80001f38
    mem[1999] <= 16'h0004; // 0x80001f3c
    mem[2000] <= 16'h0024; // 0x80001f40
    mem[2001] <= 16'h0097; // 0x80001f44
    mem[2002] <= 16'h0017; // 0x80001f48
    mem[2003] <= 16'h0014; // 0x80001f4c
    mem[2004] <= 16'h01d4; // 0x80001f50
    mem[2005] <= 16'h0007; // 0x80001f54
    mem[2006] <= 16'hfd04; // 0x80001f58
    mem[2007] <= 16'hfd0e; // 0x80001f5c
    mem[2008] <= 16'hfee5; // 0x80001f60
    mem[2009] <= 16'h000e; // 0x80001f64
    mem[2010] <= 16'hf95f; // 0x80001f68
    mem[2011] <= 16'h1a08; // 0x80001f6c
    mem[2012] <= 16'h0006; // 0x80001f70
    mem[2013] <= 16'h0009; // 0x80001f74
    mem[2014] <= 16'h0046; // 0x80001f78
    mem[2015] <= 16'h00c1; // 0x80001f7c
    mem[2016] <= 16'hdb8f; // 0x80001f80
    mem[2017] <= 16'he59f; // 0x80001f84
    mem[2018] <= 16'h1c08; // 0x80001f88
    mem[2019] <= 16'h0080; // 0x80001f8c
    mem[2020] <= 16'hf1df; // 0x80001f90
    mem[2021] <= 16'h1a08; // 0x80001f94
    mem[2022] <= 16'h000a; // 0x80001f98
    mem[2023] <= 16'h0009; // 0x80001f9c
    mem[2024] <= 16'hd98f; // 0x80001fa0
    mem[2025] <= 16'h0009; // 0x80001fa4
    mem[2026] <= 16'h0780; // 0x80001fa8
    mem[2027] <= 16'hd8cf; // 0x80001fac
    mem[2028] <= 16'h0100; // 0x80001fb0
    mem[2029] <= 16'h0010; // 0x80001fb4
    mem[2030] <= 16'hef5f; // 0x80001fb8
    mem[2031] <= 16'h1608; // 0x80001fbc
    mem[2032] <= 16'h0046; // 0x80001fc0
    mem[2033] <= 16'h00f1; // 0x80001fc4
    mem[2034] <= 16'h0006; // 0x80001fc8
    mem[2035] <= 16'h120c; // 0x80001fcc
    mem[2036] <= 16'h0580; // 0x80001fd0
    mem[2037] <= 16'h02d0; // 0x80001fd4
    mem[2038] <= 16'h10fb; // 0x80001fd8
    mem[2039] <= 16'h0004; // 0x80001fdc
    mem[2040] <= 16'h000c; // 0x80001fe0
    mem[2041] <= 16'hd6df; // 0x80001fe4
    mem[2042] <= 16'h40ac; // 0x80001fe8
    mem[2043] <= 16'h0380; // 0x80001fec
    mem[2044] <= 16'h000c; // 0x80001ff0
    mem[2045] <= 16'hfffd; // 0x80001ff4
    mem[2046] <= 16'h0009; // 0x80001ff8
    mem[2047] <= 16'h000b; // 0x80001ffc
    mem[2048] <= 16'hd38f; // 0x80002000
    mem[2049] <= 16'hfe0d; // 0x80002004
    mem[2050] <= 16'hfffc; // 0x80002008
    mem[2051] <= 16'h418b; // 0x8000200c
    mem[2052] <= 16'h00fc; // 0x80002010
    mem[2053] <= 16'h000c; // 0x80002014
    mem[2054] <= 16'hdc05; // 0x80002018
    mem[2055] <= 16'h0004; // 0x8000201c
    mem[2056] <= 16'hfff4; // 0x80002020
    mem[2057] <= 16'h0144; // 0x80002024
    mem[2058] <= 16'h0009; // 0x80002028
    mem[2059] <= 16'h001c; // 0x8000202c
    mem[2060] <= 16'hd08f; // 0x80002030
    mem[2061] <= 16'h000c; // 0x80002034
    mem[2062] <= 16'hfffc; // 0x80002038
    mem[2063] <= 16'hfe05; // 0x8000203c
    mem[2064] <= 16'hd980; // 0x80002040
    mem[2065] <= 16'h0200; // 0x80002044
    mem[2066] <= 16'hfffc; // 0x80002048
    mem[2067] <= 16'h0009; // 0x8000204c
    mem[2068] <= 16'h0004; // 0x80002050
    mem[2069] <= 16'hce4f; // 0x80002054
    mem[2070] <= 16'hfe0c; // 0x80002058
    mem[2071] <= 16'hd81f; // 0x8000205c
    mem[2072] <= 16'h0c08; // 0x80002060
    mem[2073] <= 16'h00a0; // 0x80002064
    mem[2074] <= 16'he45f; // 0x80002068
    mem[2075] <= 16'h1008; // 0x8000206c
    mem[2076] <= 16'h00c1; // 0x80002070
    mem[2077] <= 16'hc80f; // 0x80002074
    mem[2078] <= 16'h0005; // 0x80002078
    mem[2079] <= 16'h0005; // 0x8000207c
    mem[2080] <= 16'h00a0; // 0x80002080
    mem[2081] <= 16'he205; // 0x80002084
    mem[2082] <= 16'h00b1; // 0x80002088
    mem[2083] <= 16'h00a1; // 0x8000208c
    mem[2084] <= 16'h0009; // 0x80002090
    mem[2085] <= 16'h02d0; // 0x80002094
    mem[2086] <= 16'hca0f; // 0x80002098
    mem[2087] <= 16'h0041; // 0x8000209c
    mem[2088] <= 16'h0081; // 0x800020a0
    mem[2089] <= 16'h40c0; // 0x800020a4
    mem[2090] <= 16'h00c0; // 0x800020a8
    mem[2091] <= 16'h40d0; // 0x800020ac
    mem[2092] <= 16'h40f6; // 0x800020b0
    mem[2093] <= 16'he09f; // 0x800020b4
    mem[2094] <= 16'h0017; // 0x800020b8
    mem[2095] <= 16'h0015; // 0x800020bc
    mem[2096] <= 16'h0004; // 0x800020c0
    mem[2097] <= 16'hd71f; // 0x800020c4
    mem[2098] <= 16'h0808; // 0x800020c8
    mem[2099] <= 16'h0009; // 0x800020cc
    mem[2100] <= 16'h0250; // 0x800020d0
    mem[2101] <= 16'hc64f; // 0x800020d4
    mem[2102] <= 16'h000c; // 0x800020d8
    mem[2103] <= 16'hd01f; // 0x800020dc
    mem[2104] <= 16'h000c; // 0x800020e0
    mem[2105] <= 16'hf205; // 0x800020e4
    mem[2106] <= 16'hf5df; // 0x800020e8
    mem[2107] <= 16'h0380; // 0x800020ec
    mem[2108] <= 16'h02d0; // 0x800020f0
    mem[2109] <= 16'h0000; // 0x800020f4
    mem[2110] <= 16'h378c; // 0x800020f8
    mem[2111] <= 16'h0280; // 0x800020fc
    mem[2112] <= 16'hecfb; // 0x80002100
    mem[2113] <= 16'hf19f; // 0x80002104
    mem[2114] <= 16'h000e; // 0x80002108
    mem[2115] <= 16'h0004; // 0x8000210c
    mem[2116] <= 16'hdedf; // 0x80002110
    mem[2117] <= 16'h0280; // 0x80002114
    mem[2118] <= 16'h0000; // 0x80002118
    mem[2119] <= 16'h354c; // 0x8000211c
    mem[2120] <= 16'hefdf; // 0x80002120
    mem[2121] <= 16'h0008; // 0x80002124
    mem[2122] <= 16'he49f; // 0x80002128
    mem[2123] <= 16'h0111; // 0x8000212c
    mem[2124] <= 16'h00a0; // 0x80002130
    mem[2125] <= 16'hd79f; // 0x80002134
    mem[2126] <= 16'h0008; // 0x80002138
    mem[2127] <= 16'he85f; // 0x8000213c
    mem[2128] <= 16'h0111; // 0x80002140
    mem[2129] <= 16'he55f; // 0x80002144
    mem[2130] <= 16'h0111; // 0x80002148
    mem[2131] <= 16'h0080; // 0x8000214c
    mem[2132] <= 16'hd5df; // 0x80002150
    mem[2133] <= 16'h0111; // 0x80002154
    mem[2134] <= 16'hd81f; // 0x80002158
    mem[2135] <= 16'h0111; // 0x8000215c
    mem[2136] <= 16'hd49f; // 0x80002160
    mem[2137] <= 16'h0111; // 0x80002164
    mem[2138] <= 16'hf65f; // 0x80002168
    mem[2139] <= 16'h0111; // 0x8000216c
    mem[2140] <= 16'hf01f; // 0x80002170
    mem[2141] <= 16'hfb01; // 0x80002174
    mem[2142] <= 16'h0381; // 0x80002178
    mem[2143] <= 16'h0281; // 0x8000217c
    mem[2144] <= 16'h00a1; // 0x80002180
    mem[2145] <= 16'h02c1; // 0x80002184
    mem[2146] <= 16'h0005; // 0x80002188
    mem[2147] <= 16'h0003; // 0x8000218c
    mem[2148] <= 16'h00c1; // 0x80002190
    mem[2149] <= 16'h0211; // 0x80002194
    mem[2150] <= 16'h04f1; // 0x80002198
    mem[2151] <= 16'h02d1; // 0x8000219c
    mem[2152] <= 16'h04e1; // 0x800021a0
    mem[2153] <= 16'h0501; // 0x800021a4
    mem[2154] <= 16'h0511; // 0x800021a8
    mem[2155] <= 16'h0061; // 0x800021ac
    mem[2156] <= 16'hbd9f; // 0x800021b0
    mem[2157] <= 16'h00c1; // 0x800021b4
    mem[2158] <= 16'h0007; // 0x800021b8
    mem[2159] <= 16'h00c1; // 0x800021bc
    mem[2160] <= 16'h02c1; // 0x800021c0
    mem[2161] <= 16'h4085; // 0x800021c4
    mem[2162] <= 16'h0281; // 0x800021c8
    mem[2163] <= 16'h0501; // 0x800021cc
    mem[2164] <= 16'h0000; // 0x800021d0
    mem[2165] <= 16'hfe01; // 0x800021d4
    mem[2166] <= 16'h0011; // 0x800021d8
    mem[2167] <= 16'h0081; // 0x800021dc
    mem[2168] <= 16'h0091; // 0x800021e0
    mem[2169] <= 16'h0201; // 0x800021e4
    mem[2170] <= 16'h0121; // 0x800021e8
    mem[2171] <= 16'h0131; // 0x800021ec
    mem[2172] <= 16'hf801; // 0x800021f0
    mem[2173] <= 16'h0005; // 0x800021f4
    mem[2174] <= 16'h0005; // 0x800021f8
    mem[2175] <= 16'h841f; // 0x800021fc
    mem[2176] <= 16'h0009; // 0x80002200
    mem[2177] <= 16'h0009; // 0x80002204
    mem[2178] <= 16'hea0f; // 0x80002208
    mem[2179] <= 16'h0000; // 0x8000220c
    mem[2180] <= 16'h0000; // 0x80002210
    mem[2181] <= 16'h6310; // 0x80002214
    mem[2182] <= 16'h03f1; // 0x80002218
    mem[2183] <= 16'h0000; // 0x8000221c
    mem[2184] <= 16'h2e46; // 0x80002220
    mem[2185] <= 16'hfc04; // 0x80002224
    mem[2186] <= 16'h0005; // 0x80002228
    mem[2187] <= 16'h0406; // 0x8000222c
    mem[2188] <= 16'h0000; // 0x80002230
    mem[2189] <= 16'h2d46; // 0x80002234
    mem[2190] <= 16'h0004; // 0x80002238
    mem[2191] <= 16'h0206; // 0x8000223c
    mem[2192] <= 16'h0009; // 0x80002240
    mem[2193] <= 16'h0000; // 0x80002244
    mem[2194] <= 16'h2b86; // 0x80002248
    mem[2195] <= 16'h0000; // 0x8000224c
    mem[2196] <= 16'h2285; // 0x80002250
    mem[2197] <= 16'hf21f; // 0x80002254
    mem[2198] <= 16'h00a9; // 0x80002258
    mem[2199] <= 16'h0124; // 0x8000225c
    mem[2200] <= 16'h0004; // 0x80002260
    mem[2201] <= 16'h861f; // 0x80002264
    mem[2202] <= 16'h0009; // 0x80002268
    mem[2203] <= 16'he20f; // 0x8000226c
    mem[2204] <= 16'h0000; // 0x80002270
    mem[2205] <= 16'h2886; // 0x80002274
    mem[2206] <= 16'h0000; // 0x80002278
    mem[2207] <= 16'h1fc5; // 0x8000227c
    mem[2208] <= 16'h0004; // 0x80002280
    mem[2209] <= 16'hef1f; // 0x80002284
    mem[2210] <= 16'h0000; // 0x80002288
    mem[2211] <= 16'h27c6; // 0x8000228c
    mem[2212] <= 16'h00a4; // 0x80002290
    mem[2213] <= 16'hfc06; // 0x80002294
    mem[2214] <= 16'hfa9f; // 0x80002298
    mem[2215] <= 16'hfc01; // 0x8000229c
    mem[2216] <= 16'h0281; // 0x800022a0
    mem[2217] <= 16'h0321; // 0x800022a4
    mem[2218] <= 16'h0331; // 0x800022a8
    mem[2219] <= 16'h0341; // 0x800022ac
    mem[2220] <= 16'h0351; // 0x800022b0
    mem[2221] <= 16'h0211; // 0x800022b4
    mem[2222] <= 16'h0291; // 0x800022b8
    mem[2223] <= 16'h0361; // 0x800022bc
    mem[2224] <= 16'h0171; // 0x800022c0
    mem[2225] <= 16'h0181; // 0x800022c4
    mem[2226] <= 16'h0191; // 0x800022c8
    mem[2227] <= 16'h0005; // 0x800022cc
    mem[2228] <= 16'h00b1; // 0x800022d0
    mem[2229] <= 16'h0000; // 0x800022d4
    mem[2230] <= 16'hf149; // 0x800022d8
    mem[2231] <= 16'h0010; // 0x800022dc
    mem[2232] <= 16'h0300; // 0x800022e0
    mem[2233] <= 16'hfff0; // 0x800022e4
    mem[2234] <= 16'h0004; // 0x800022e8
    mem[2235] <= 16'h0250; // 0x800022ec
    mem[2236] <= 16'h0095; // 0x800022f0
    mem[2237] <= 16'h0605; // 0x800022f4
    mem[2238] <= 16'h0000; // 0x800022f8
    mem[2239] <= 16'h0014; // 0x800022fc
    mem[2240] <= 16'h970f; // 0x80002300
    mem[2241] <= 16'h0004; // 0x80002304
    mem[2242] <= 16'hfe95; // 0x80002308
    mem[2243] <= 16'h00c1; // 0x8000230c
    mem[2244] <= 16'h0014; // 0x80002310
    mem[2245] <= 16'h0014; // 0x80002314
    mem[2246] <= 16'hfff0; // 0x80002318
    mem[2247] <= 16'h0006; // 0x8000231c
    mem[2248] <= 16'h000c; // 0x80002320
    mem[2249] <= 16'h0000; // 0x80002324
    mem[2250] <= 16'h0200; // 0x80002328
    mem[2251] <= 16'h0004; // 0x8000232c
    mem[2252] <= 16'h0000; // 0x80002330
    mem[2253] <= 16'h0550; // 0x80002334
    mem[2254] <= 16'h0090; // 0x80002338
    mem[2255] <= 16'h02d0; // 0x8000233c
    mem[2256] <= 16'hfdde; // 0x80002340
    mem[2257] <= 16'h0ff7; // 0x80002344
    mem[2258] <= 16'h0017; // 0x80002348
    mem[2259] <= 16'h26f6; // 0x8000234c
    mem[2260] <= 16'h0027; // 0x80002350
    mem[2261] <= 16'h0127; // 0x80002354
    mem[2262] <= 16'h0007; // 0x80002358
    mem[2263] <= 16'h0127; // 0x8000235c
    mem[2264] <= 16'h0007; // 0x80002360
    mem[2265] <= 16'h03c1; // 0x80002364
    mem[2266] <= 16'h0381; // 0x80002368
    mem[2267] <= 16'h0341; // 0x8000236c
    mem[2268] <= 16'h0301; // 0x80002370
    mem[2269] <= 16'h02c1; // 0x80002374
    mem[2270] <= 16'h0281; // 0x80002378
    mem[2271] <= 16'h0241; // 0x8000237c
    mem[2272] <= 16'h0201; // 0x80002380
    mem[2273] <= 16'h01c1; // 0x80002384
    mem[2274] <= 16'h0181; // 0x80002388
    mem[2275] <= 16'h0141; // 0x8000238c
    mem[2276] <= 16'h0401; // 0x80002390
    mem[2277] <= 16'h0000; // 0x80002394
    mem[2278] <= 16'h000b; // 0x80002398
    mem[2279] <= 16'h0000; // 0x8000239c
    mem[2280] <= 16'h0017; // 0x800023a0
    mem[2281] <= 16'h0004; // 0x800023a4
    mem[2282] <= 16'hf99f; // 0x800023a8
    mem[2283] <= 16'h2a08; // 0x800023ac
    mem[2284] <= 16'h0100; // 0x800023b0
    mem[2285] <= 16'h00c1; // 0x800023b4
    mem[2286] <= 16'h8e0f; // 0x800023b8
    mem[2287] <= 16'h0005; // 0x800023bc
    mem[2288] <= 16'h0005; // 0x800023c0
    mem[2289] <= 16'h000b; // 0x800023c4
    mem[2290] <= 16'h000b; // 0x800023c8
    mem[2291] <= 16'h000c; // 0x800023cc
    mem[2292] <= 16'h000c; // 0x800023d0
    mem[2293] <= 16'h0004; // 0x800023d4
    mem[2294] <= 16'h978f; // 0x800023d8
    mem[2295] <= 16'hf0df; // 0x800023dc
    mem[2296] <= 16'h2608; // 0x800023e0
    mem[2297] <= 16'h0000; // 0x800023e4
    mem[2298] <= 16'h0250; // 0x800023e8
    mem[2299] <= 16'h884f; // 0x800023ec
    mem[2300] <= 16'hef9f; // 0x800023f0
    mem[2301] <= 16'h0008; // 0x800023f4
    mem[2302] <= 16'h0017; // 0x800023f8
    mem[2303] <= 16'h0048; // 0x800023fc
    mem[2304] <= 16'h0004; // 0x80002400
    mem[2305] <= 16'h000a; // 0x80002404
    mem[2306] <= 16'hf20b; // 0x80002408
    mem[2307] <= 16'h0004; // 0x8000240c
    mem[2308] <= 16'hfff0; // 0x80002410
    mem[2309] <= 16'hf2df; // 0x80002414
    mem[2310] <= 16'h0017; // 0x80002418
    mem[2311] <= 16'h0003; // 0x8000241c
    mem[2312] <= 16'h0004; // 0x80002420
    mem[2313] <= 16'hf1df; // 0x80002424
    mem[2314] <= 16'h0017; // 0x80002428
    mem[2315] <= 16'h000a; // 0x8000242c
    mem[2316] <= 16'h0004; // 0x80002430
    mem[2317] <= 16'hf0df; // 0x80002434
    mem[2318] <= 16'h0017; // 0x80002438
    mem[2319] <= 16'hfd0e; // 0x8000243c
    mem[2320] <= 16'hfd0e; // 0x80002440
    mem[2321] <= 16'h1cf5; // 0x80002444
    mem[2322] <= 16'h0004; // 0x80002448
    mem[2323] <= 16'h0024; // 0x8000244c
    mem[2324] <= 16'h0097; // 0x80002450
    mem[2325] <= 16'h0017; // 0x80002454
    mem[2326] <= 16'h0014; // 0x80002458
    mem[2327] <= 16'h01d4; // 0x8000245c
    mem[2328] <= 16'h0007; // 0x80002460
    mem[2329] <= 16'hfd04; // 0x80002464
    mem[2330] <= 16'hfd0e; // 0x80002468
    mem[2331] <= 16'hfef5; // 0x8000246c
    mem[2332] <= 16'h000e; // 0x80002470
    mem[2333] <= 16'hf95f; // 0x80002474
    mem[2334] <= 16'h1a08; // 0x80002478
    mem[2335] <= 16'h0006; // 0x8000247c
    mem[2336] <= 16'h0000; // 0x80002480
    mem[2337] <= 16'h0046; // 0x80002484
    mem[2338] <= 16'h00c1; // 0x80002488
    mem[2339] <= 16'hfe5f; // 0x8000248c
    mem[2340] <= 16'he59f; // 0x80002490
    mem[2341] <= 16'h1a08; // 0x80002494
    mem[2342] <= 16'h0080; // 0x80002498
    mem[2343] <= 16'hf19f; // 0x8000249c
    mem[2344] <= 16'h1808; // 0x800024a0
    mem[2345] <= 16'h0000; // 0x800024a4
    mem[2346] <= 16'h000a; // 0x800024a8
    mem[2347] <= 16'hfc5f; // 0x800024ac
    mem[2348] <= 16'h0000; // 0x800024b0
    mem[2349] <= 16'h0780; // 0x800024b4
    mem[2350] <= 16'hfb9f; // 0x800024b8
    mem[2351] <= 16'h0100; // 0x800024bc
    mem[2352] <= 16'h0010; // 0x800024c0
    mem[2353] <= 16'hef1f; // 0x800024c4
    mem[2354] <= 16'h1608; // 0x800024c8
    mem[2355] <= 16'h0046; // 0x800024cc
    mem[2356] <= 16'h00f1; // 0x800024d0
    mem[2357] <= 16'h0006; // 0x800024d4
    mem[2358] <= 16'h100c; // 0x800024d8
    mem[2359] <= 16'h0570; // 0x800024dc
    mem[2360] <= 16'h02d0; // 0x800024e0
    mem[2361] <= 16'h0efb; // 0x800024e4
    mem[2362] <= 16'h0004; // 0x800024e8
    mem[2363] <= 16'h000c; // 0x800024ec
    mem[2364] <= 16'h861f; // 0x800024f0
    mem[2365] <= 16'h40ab; // 0x800024f4
    mem[2366] <= 16'h0370; // 0x800024f8
    mem[2367] <= 16'h000b; // 0x800024fc
    mem[2368] <= 16'hfffc; // 0x80002500
    mem[2369] <= 16'h0000; // 0x80002504
    mem[2370] <= 16'h000b; // 0x80002508
    mem[2371] <= 16'hf65f; // 0x8000250c
    mem[2372] <= 16'hfe0c; // 0x80002510
    mem[2373] <= 16'hfffb; // 0x80002514
    mem[2374] <= 16'h417a; // 0x80002518
    mem[2375] <= 16'h00fb; // 0x8000251c
    mem[2376] <= 16'h000c; // 0x80002520
    mem[2377] <= 16'hdc05; // 0x80002524
    mem[2378] <= 16'h0004; // 0x80002528
    mem[2379] <= 16'hfff4; // 0x8000252c
    mem[2380] <= 16'h0134; // 0x80002530
    mem[2381] <= 16'h0000; // 0x80002534
    mem[2382] <= 16'h001c; // 0x80002538
    mem[2383] <= 16'hf35f; // 0x8000253c
    mem[2384] <= 16'h000c; // 0x80002540
    mem[2385] <= 16'hfffb; // 0x80002544
    mem[2386] <= 16'hfe05; // 0x80002548
    mem[2387] <= 16'hd970; // 0x8000254c
    mem[2388] <= 16'h0200; // 0x80002550
    mem[2389] <= 16'hfffb; // 0x80002554
    mem[2390] <= 16'h0000; // 0x80002558
    mem[2391] <= 16'h0004; // 0x8000255c
    mem[2392] <= 16'hf11f; // 0x80002560
    mem[2393] <= 16'hfe0b; // 0x80002564
    mem[2394] <= 16'hd81f; // 0x80002568
    mem[2395] <= 16'h0a08; // 0x8000256c
    mem[2396] <= 16'h00a0; // 0x80002570
    mem[2397] <= 16'he41f; // 0x80002574
    mem[2398] <= 16'h0e08; // 0x80002578
    mem[2399] <= 16'h00c1; // 0x8000257c
    mem[2400] <= 16'hf75f; // 0x80002580
    mem[2401] <= 16'h0005; // 0x80002584
    mem[2402] <= 16'h0005; // 0x80002588
    mem[2403] <= 16'h00a0; // 0x8000258c
    mem[2404] <= 16'he205; // 0x80002590
    mem[2405] <= 16'h0000; // 0x80002594
    mem[2406] <= 16'h02d0; // 0x80002598
    mem[2407] <= 16'hed5f; // 0x8000259c
    mem[2408] <= 16'h4180; // 0x800025a0
    mem[2409] <= 16'h0180; // 0x800025a4
    mem[2410] <= 16'h4090; // 0x800025a8
    mem[2411] <= 16'h40f4; // 0x800025ac
    mem[2412] <= 16'he15f; // 0x800025b0
    mem[2413] <= 16'h0017; // 0x800025b4
    mem[2414] <= 16'h0015; // 0x800025b8
    mem[2415] <= 16'h0004; // 0x800025bc
    mem[2416] <= 16'hd81f; // 0x800025c0
    mem[2417] <= 16'h0808; // 0x800025c4
    mem[2418] <= 16'h0000; // 0x800025c8
    mem[2419] <= 16'h0250; // 0x800025cc
    mem[2420] <= 16'hea1f; // 0x800025d0
    mem[2421] <= 16'h000c; // 0x800025d4
    mem[2422] <= 16'hd11f; // 0x800025d8
    mem[2423] <= 16'h000c; // 0x800025dc
    mem[2424] <= 16'hf405; // 0x800025e0
    mem[2425] <= 16'hf6df; // 0x800025e4
    mem[2426] <= 16'h0370; // 0x800025e8
    mem[2427] <= 16'h02d0; // 0x800025ec
    mem[2428] <= 16'h0000; // 0x800025f0
    mem[2429] <= 16'he7cc; // 0x800025f4
    mem[2430] <= 16'h0280; // 0x800025f8
    mem[2431] <= 16'heefb; // 0x800025fc
    mem[2432] <= 16'hf29f; // 0x80002600
    mem[2433] <= 16'h000e; // 0x80002604
    mem[2434] <= 16'h0004; // 0x80002608
    mem[2435] <= 16'hdfdf; // 0x8000260c
    mem[2436] <= 16'h0280; // 0x80002610
    mem[2437] <= 16'h0000; // 0x80002614
    mem[2438] <= 16'he58c; // 0x80002618
    mem[2439] <= 16'hf0df; // 0x8000261c
    mem[2440] <= 16'h0008; // 0x80002620
    mem[2441] <= 16'he59f; // 0x80002624
    mem[2442] <= 16'h0111; // 0x80002628
    mem[2443] <= 16'h00a0; // 0x8000262c
    mem[2444] <= 16'hd85f; // 0x80002630
    mem[2445] <= 16'h0008; // 0x80002634
    mem[2446] <= 16'he95f; // 0x80002638
    mem[2447] <= 16'h0111; // 0x8000263c
    mem[2448] <= 16'he65f; // 0x80002640
    mem[2449] <= 16'h0111; // 0x80002644
    mem[2450] <= 16'h0080; // 0x80002648
    mem[2451] <= 16'hd69f; // 0x8000264c
    mem[2452] <= 16'h0111; // 0x80002650
    mem[2453] <= 16'hd91f; // 0x80002654
    mem[2454] <= 16'h0111; // 0x80002658
    mem[2455] <= 16'hd55f; // 0x8000265c
    mem[2456] <= 16'h0111; // 0x80002660
    mem[2457] <= 16'hf65f; // 0x80002664
    mem[2458] <= 16'h0111; // 0x80002668
    mem[2459] <= 16'hf11f; // 0x8000266c
    mem[2460] <= 16'hfc01; // 0x80002670
    mem[2461] <= 16'h0241; // 0x80002674
    mem[2462] <= 16'h02b1; // 0x80002678
    mem[2463] <= 16'h0003; // 0x8000267c
    mem[2464] <= 16'h0011; // 0x80002680
    mem[2465] <= 16'h02c1; // 0x80002684
    mem[2466] <= 16'h02d1; // 0x80002688
    mem[2467] <= 16'h02e1; // 0x8000268c
    mem[2468] <= 16'h02f1; // 0x80002690
    mem[2469] <= 16'h0301; // 0x80002694
    mem[2470] <= 16'h0311; // 0x80002698
    mem[2471] <= 16'h0061; // 0x8000269c
    mem[2472] <= 16'hbfdf; // 0x800026a0
    mem[2473] <= 16'h01c1; // 0x800026a4
    mem[2474] <= 16'h0000; // 0x800026a8
    mem[2475] <= 16'h0401; // 0x800026ac
    mem[2476] <= 16'h0000; // 0x800026b0
    mem[2477] <= 16'h0015; // 0x800026b4
    mem[2478] <= 16'hfff5; // 0x800026b8
    mem[2479] <= 16'h0015; // 0x800026bc
    mem[2480] <= 16'hfff5; // 0x800026c0
    mem[2481] <= 16'h0007; // 0x800026c4
    mem[2482] <= 16'hfee7; // 0x800026c8
    mem[2483] <= 16'h40e7; // 0x800026cc
    mem[2484] <= 16'h0000; // 0x800026d0
    mem[2485] <= 16'h0000; // 0x800026d4
    mem[2486] <= 16'hff5f; // 0x800026d8
    mem[2487] <= 16'h0005; // 0x800026dc
    mem[2488] <= 16'h0015; // 0x800026e0
    mem[2489] <= 16'hfff5; // 0x800026e4
    mem[2490] <= 16'h0017; // 0x800026e8
    mem[2491] <= 16'hfee7; // 0x800026ec
    mem[2492] <= 16'hfe07; // 0x800026f0
    mem[2493] <= 16'h0000; // 0x800026f4
    mem[2494] <= 16'h0005; // 0x800026f8
    mem[2495] <= 16'h0200; // 0x800026fc
    mem[2496] <= 16'h0005; // 0x80002700
    mem[2497] <= 16'h00d7; // 0x80002704
    mem[2498] <= 16'h0007; // 0x80002708
    mem[2499] <= 16'h0017; // 0x8000270c
    mem[2500] <= 16'h0007; // 0x80002710
    mem[2501] <= 16'hfed7; // 0x80002714
    mem[2502] <= 16'hfd57; // 0x80002718
    mem[2503] <= 16'h0fd6; // 0x8000271c
    mem[2504] <= 16'h0406; // 0x80002720
    mem[2505] <= 16'h0000; // 0x80002724
    mem[2506] <= 16'h0407; // 0x80002728
    mem[2507] <= 16'h0000; // 0x8000272c
    mem[2508] <= 16'h0017; // 0x80002730
    mem[2509] <= 16'h0026; // 0x80002734
    mem[2510] <= 16'hfd07; // 0x80002738
    mem[2511] <= 16'h0007; // 0x8000273c
    mem[2512] <= 16'h00d5; // 0x80002740
    mem[2513] <= 16'h0015; // 0x80002744
    mem[2514] <= 16'h00a6; // 0x80002748
    mem[2515] <= 16'hfe07; // 0x8000274c
    mem[2516] <= 16'h0005; // 0x80002750
    mem[2517] <= 16'h40d0; // 0x80002754
    mem[2518] <= 16'h0006; // 0x80002758
    mem[2519] <= 16'h0000; // 0x8000275c
    mem[2520] <= 16'hfd37; // 0x80002760
    mem[2521] <= 16'h0017; // 0x80002764
    mem[2522] <= 16'h0015; // 0x80002768
    mem[2523] <= 16'h0017; // 0x8000276c
    mem[2524] <= 16'hfa07; // 0x80002770
    mem[2525] <= 16'h0000; // 0x80002774
    mem[2526] <= 16'hfd9f; // 0x80002778
    mem[2527] <= 16'h0000; // 0x8000277c
    mem[2528] <= 16'hfd9f; // 0x80002780
    mem[2529] <= 16'h0006; // 0x80002784
    mem[2530] <= 16'h0006; // 0x80002788
    mem[2531] <= 16'h0005; // 0x8000278c
    mem[2532] <= 16'h0005; // 0x80002790
    mem[2533] <= 16'h0c06; // 0x80002794
    mem[2534] <= 16'h12c5; // 0x80002798
    mem[2535] <= 16'h0001; // 0x8000279c
    mem[2536] <= 16'h22f6; // 0x800027a0
    mem[2537] <= 16'h0ff0; // 0x800027a4
    mem[2538] <= 16'h00c7; // 0x800027a8
    mem[2539] <= 16'h0080; // 0x800027ac
    mem[2540] <= 16'h8000; // 0x800027b0
    mem[2541] <= 16'h0066; // 0x800027b4
    mem[2542] <= 16'h3407; // 0x800027b8
    mem[2543] <= 16'h00e7; // 0x800027bc
    mem[2544] <= 16'h0007; // 0x800027c0
    mem[2545] <= 16'h0067; // 0x800027c4
    mem[2546] <= 16'h0200; // 0x800027c8
    mem[2547] <= 16'h4067; // 0x800027cc
    mem[2548] <= 16'h0007; // 0x800027d0
    mem[2549] <= 16'h00f5; // 0x800027d4
    mem[2550] <= 16'h0065; // 0x800027d8
    mem[2551] <= 16'h00f6; // 0x800027dc
    mem[2552] <= 16'h00e3; // 0x800027e0
    mem[2553] <= 16'h00f5; // 0x800027e4
    mem[2554] <= 16'h0108; // 0x800027e8
    mem[2555] <= 16'h02b8; // 0x800027ec
    mem[2556] <= 16'h0108; // 0x800027f0
    mem[2557] <= 16'h0106; // 0x800027f4
    mem[2558] <= 16'h010e; // 0x800027f8
    mem[2559] <= 16'h02b8; // 0x800027fc
    mem[2560] <= 16'h02e6; // 0x80002800
    mem[2561] <= 16'h0106; // 0x80002804
    mem[2562] <= 16'h00f6; // 0x80002808
    mem[2563] <= 16'h00a8; // 0x8000280c
    mem[2564] <= 16'h0118; // 0x80002810
    mem[2565] <= 16'hfff7; // 0x80002814
    mem[2566] <= 16'h0118; // 0x80002818
    mem[2567] <= 16'h3ca8; // 0x8000281c
    mem[2568] <= 16'h0007; // 0x80002820
    mem[2569] <= 16'h40a8; // 0x80002824
    mem[2570] <= 16'h02b8; // 0x80002828
    mem[2571] <= 16'h010e; // 0x8000282c
    mem[2572] <= 16'h010e; // 0x80002830
    mem[2573] <= 16'h02b8; // 0x80002834
    mem[2574] <= 16'h02a6; // 0x80002838
    mem[2575] <= 16'h0108; // 0x8000283c
    mem[2576] <= 16'h01c8; // 0x80002840
    mem[2577] <= 16'h00c8; // 0x80002844
    mem[2578] <= 16'h0108; // 0x80002848
    mem[2579] <= 16'hfff5; // 0x8000284c
    mem[2580] <= 16'h3318; // 0x80002850
    mem[2581] <= 16'hffe5; // 0x80002854
    mem[2582] <= 16'h32c8; // 0x80002858
    mem[2583] <= 16'h0107; // 0x8000285c
    mem[2584] <= 16'h00a7; // 0x80002860
    mem[2585] <= 16'h0000; // 0x80002864
    mem[2586] <= 16'h0007; // 0x80002868
    mem[2587] <= 16'h0000; // 0x8000286c
    mem[2588] <= 16'h12d5; // 0x80002870
    mem[2589] <= 16'h0001; // 0x80002874
    mem[2590] <= 16'h12f6; // 0x80002878
    mem[2591] <= 16'h0100; // 0x8000287c
    mem[2592] <= 16'h0180; // 0x80002880
    mem[2593] <= 16'h00e6; // 0x80002884
    mem[2594] <= 16'h0100; // 0x80002888
    mem[2595] <= 16'h8000; // 0x8000288c
    mem[2596] <= 16'h00f6; // 0x80002890
    mem[2597] <= 16'h3408; // 0x80002894
    mem[2598] <= 16'h0117; // 0x80002898
    mem[2599] <= 16'h0007; // 0x8000289c
    mem[2600] <= 16'h0200; // 0x800028a0
    mem[2601] <= 16'h00fe; // 0x800028a4
    mem[2602] <= 16'h41ce; // 0x800028a8
    mem[2603] <= 16'h120e; // 0x800028ac
    mem[2604] <= 16'h0000; // 0x800028b0
    mem[2605] <= 16'h0010; // 0x800028b4
    mem[2606] <= 16'h0f03; // 0x800028b8
    mem[2607] <= 16'h00c5; // 0x800028bc
    mem[2608] <= 16'h0017; // 0x800028c0
    mem[2609] <= 16'h0e00; // 0x800028c4
    mem[2610] <= 16'h0006; // 0x800028c8
    mem[2611] <= 16'h0010; // 0x800028cc
    mem[2612] <= 16'h02c8; // 0x800028d0
    mem[2613] <= 16'h0001; // 0x800028d4
    mem[2614] <= 16'h0ef8; // 0x800028d8
    mem[2615] <= 16'h0100; // 0x800028dc
    mem[2616] <= 16'h0180; // 0x800028e0
    mem[2617] <= 16'h00f8; // 0x800028e4
    mem[2618] <= 16'h0100; // 0x800028e8
    mem[2619] <= 16'h8000; // 0x800028ec
    mem[2620] <= 16'h0068; // 0x800028f0
    mem[2621] <= 16'h3407; // 0x800028f4
    mem[2622] <= 16'h00e7; // 0x800028f8
    mem[2623] <= 16'h0007; // 0x800028fc
    mem[2624] <= 16'h0067; // 0x80002900
    mem[2625] <= 16'h0200; // 0x80002904
    mem[2626] <= 16'h4067; // 0x80002908
    mem[2627] <= 16'h1c07; // 0x8000290c
    mem[2628] <= 16'h0108; // 0x80002910
    mem[2629] <= 16'h4115; // 0x80002914
    mem[2630] <= 16'h0108; // 0x80002918
    mem[2631] <= 16'h010f; // 0x8000291c
    mem[2632] <= 16'h0010; // 0x80002920
    mem[2633] <= 16'h010e; // 0x80002924
    mem[2634] <= 16'h03d7; // 0x80002928
    mem[2635] <= 16'h03d7; // 0x8000292c
    mem[2636] <= 16'h03e6; // 0x80002930
    mem[2637] <= 16'h0107; // 0x80002934
    mem[2638] <= 16'h00f7; // 0x80002938
    mem[2639] <= 16'h00c7; // 0x8000293c
    mem[2640] <= 16'h0117; // 0x80002940
    mem[2641] <= 16'hfff6; // 0x80002944
    mem[2642] <= 16'h0117; // 0x80002948
    mem[2643] <= 16'h28c7; // 0x8000294c
    mem[2644] <= 16'h0007; // 0x80002950
    mem[2645] <= 16'h40c7; // 0x80002954
    mem[2646] <= 16'h03d7; // 0x80002958
    mem[2647] <= 16'h010e; // 0x8000295c
    mem[2648] <= 16'h010e; // 0x80002960
    mem[2649] <= 16'h03d7; // 0x80002964
    mem[2650] <= 16'h03e5; // 0x80002968
    mem[2651] <= 16'h0107; // 0x8000296c
    mem[2652] <= 16'h01c7; // 0x80002970
    mem[2653] <= 16'h01e7; // 0x80002974
    mem[2654] <= 16'h00f8; // 0x80002978
    mem[2655] <= 16'hfff5; // 0x8000297c
    mem[2656] <= 16'h1f17; // 0x80002980
    mem[2657] <= 16'hffe5; // 0x80002984
    mem[2658] <= 16'h1fe7; // 0x80002988
    mem[2659] <= 16'h0106; // 0x8000298c
    mem[2660] <= 16'h00a7; // 0x80002990
    mem[2661] <= 16'h0007; // 0x80002994
    mem[2662] <= 16'h0000; // 0x80002998
    mem[2663] <= 16'h0000; // 0x8000299c
    mem[2664] <= 16'h0000; // 0x800029a0
    mem[2665] <= 16'h0007; // 0x800029a4
    mem[2666] <= 16'h0000; // 0x800029a8
    mem[2667] <= 16'h0ff0; // 0x800029ac
    mem[2668] <= 16'h00de; // 0x800029b0
    mem[2669] <= 16'h0037; // 0x800029b4
    mem[2670] <= 16'hed5f; // 0x800029b8
    mem[2671] <= 16'h0ff0; // 0x800029bc
    mem[2672] <= 16'hf317; // 0x800029c0
    mem[2673] <= 16'h0080; // 0x800029c4
    mem[2674] <= 16'hf25f; // 0x800029c8
    mem[2675] <= 16'h0100; // 0x800029cc
    mem[2676] <= 16'h0180; // 0x800029d0
    mem[2677] <= 16'hdcf6; // 0x800029d4
    mem[2678] <= 16'h0100; // 0x800029d8
    mem[2679] <= 16'hdd5f; // 0x800029dc
    mem[2680] <= 16'h01c6; // 0x800029e0
    mem[2681] <= 16'h01d6; // 0x800029e4
    mem[2682] <= 16'h00d8; // 0x800029e8
    mem[2683] <= 16'h01c5; // 0x800029ec
    mem[2684] <= 16'h0108; // 0x800029f0
    mem[2685] <= 16'h03e8; // 0x800029f4
    mem[2686] <= 16'h0108; // 0x800029f8
    mem[2687] <= 16'h0107; // 0x800029fc
    mem[2688] <= 16'h01d5; // 0x80002a00
    mem[2689] <= 16'h01c5; // 0x80002a04
    mem[2690] <= 16'h00be; // 0x80002a08
    mem[2691] <= 16'h0105; // 0x80002a0c
    mem[2692] <= 16'h01d6; // 0x80002a10
    mem[2693] <= 16'h03e8; // 0x80002a14
    mem[2694] <= 16'h0267; // 0x80002a18
    mem[2695] <= 16'h0108; // 0x80002a1c
    mem[2696] <= 16'h00d8; // 0x80002a20
    mem[2697] <= 16'h00f6; // 0x80002a24
    mem[2698] <= 16'h0106; // 0x80002a28
    mem[2699] <= 16'hfff3; // 0x80002a2c
    mem[2700] <= 16'h1906; // 0x80002a30
    mem[2701] <= 16'h0008; // 0x80002a34
    mem[2702] <= 16'h40f6; // 0x80002a38
    mem[2703] <= 16'h03e6; // 0x80002a3c
    mem[2704] <= 16'h0105; // 0x80002a40
    mem[2705] <= 16'h0105; // 0x80002a44
    mem[2706] <= 16'h03e6; // 0x80002a48
    mem[2707] <= 16'h03c7; // 0x80002a4c
    mem[2708] <= 16'h0106; // 0x80002a50
    mem[2709] <= 16'h00b6; // 0x80002a54
    mem[2710] <= 16'h0117; // 0x80002a58
    mem[2711] <= 16'h0107; // 0x80002a5c
    mem[2712] <= 16'hfffe; // 0x80002a60
    mem[2713] <= 16'h1507; // 0x80002a64
    mem[2714] <= 16'h0007; // 0x80002a68
    mem[2715] <= 16'h0103; // 0x80002a6c
    mem[2716] <= 16'h0001; // 0x80002a70
    mem[2717] <= 16'h01c7; // 0x80002a74
    mem[2718] <= 16'hffff; // 0x80002a78
    mem[2719] <= 16'h00d7; // 0x80002a7c
    mem[2720] <= 16'h0107; // 0x80002a80
    mem[2721] <= 16'h00d6; // 0x80002a84
    mem[2722] <= 16'h0106; // 0x80002a88
    mem[2723] <= 16'h02d5; // 0x80002a8c
    mem[2724] <= 16'h4117; // 0x80002a90
    mem[2725] <= 16'h02c5; // 0x80002a94
    mem[2726] <= 16'h010e; // 0x80002a98
    mem[2727] <= 16'h02d3; // 0x80002a9c
    mem[2728] <= 16'h00d5; // 0x80002aa0
    mem[2729] <= 16'h00b8; // 0x80002aa4
    mem[2730] <= 16'h02c3; // 0x80002aa8
    mem[2731] <= 16'h00d5; // 0x80002aac
    mem[2732] <= 16'h01e6; // 0x80002ab0
    mem[2733] <= 16'h0105; // 0x80002ab4
    mem[2734] <= 16'h00c6; // 0x80002ab8
    mem[2735] <= 16'h0ec7; // 0x80002abc
    mem[2736] <= 16'h0cc7; // 0x80002ac0
    mem[2737] <= 16'h0000; // 0x80002ac4
    mem[2738] <= 16'h0007; // 0x80002ac8
    mem[2739] <= 16'h0000; // 0x80002acc
    mem[2740] <= 16'h00f8; // 0x80002ad0
    mem[2741] <= 16'h0065; // 0x80002ad4
    mem[2742] <= 16'h0108; // 0x80002ad8
    mem[2743] <= 16'h03d6; // 0x80002adc
    mem[2744] <= 16'h0108; // 0x80002ae0
    mem[2745] <= 16'h010f; // 0x80002ae4
    mem[2746] <= 16'h00f5; // 0x80002ae8
    mem[2747] <= 16'h00f5; // 0x80002aec
    mem[2748] <= 16'h0065; // 0x80002af0
    mem[2749] <= 16'h00e3; // 0x80002af4
    mem[2750] <= 16'h0107; // 0x80002af8
    mem[2751] <= 16'h03d6; // 0x80002afc
    mem[2752] <= 16'h03ff; // 0x80002b00
    mem[2753] <= 16'h0106; // 0x80002b04
    mem[2754] <= 16'h00b6; // 0x80002b08
    mem[2755] <= 16'h00f6; // 0x80002b0c
    mem[2756] <= 16'h0116; // 0x80002b10
    mem[2757] <= 16'hffff; // 0x80002b14
    mem[2758] <= 16'h0d16; // 0x80002b18
    mem[2759] <= 16'h0af6; // 0x80002b1c
    mem[2760] <= 16'hffef; // 0x80002b20
    mem[2761] <= 16'h0116; // 0x80002b24
    mem[2762] <= 16'h40f6; // 0x80002b28
    mem[2763] <= 16'h03d6; // 0x80002b2c
    mem[2764] <= 16'h0107; // 0x80002b30
    mem[2765] <= 16'h0103; // 0x80002b34
    mem[2766] <= 16'h03d6; // 0x80002b38
    mem[2767] <= 16'h02ff; // 0x80002b3c
    mem[2768] <= 16'h0106; // 0x80002b40
    mem[2769] <= 16'h0067; // 0x80002b44
    mem[2770] <= 16'h00c7; // 0x80002b48
    mem[2771] <= 16'h0117; // 0x80002b4c
    mem[2772] <= 16'hfff7; // 0x80002b50
    mem[2773] <= 16'h0717; // 0x80002b54
    mem[2774] <= 16'h06c7; // 0x80002b58
    mem[2775] <= 16'hffe7; // 0x80002b5c
    mem[2776] <= 16'h0117; // 0x80002b60
    mem[2777] <= 16'h010f; // 0x80002b64
    mem[2778] <= 16'h40c7; // 0x80002b68
    mem[2779] <= 16'h00f5; // 0x80002b6c
    mem[2780] <= 16'hdb5f; // 0x80002b70
    mem[2781] <= 16'h0007; // 0x80002b74
    mem[2782] <= 16'he15f; // 0x80002b78
    mem[2783] <= 16'h0007; // 0x80002b7c
    mem[2784] <= 16'hcddf; // 0x80002b80
    mem[2785] <= 16'h0001; // 0x80002b84
    mem[2786] <= 16'hfff6; // 0x80002b88
    mem[2787] <= 16'h00d5; // 0x80002b8c
    mem[2788] <= 16'h0107; // 0x80002b90
    mem[2789] <= 16'h00de; // 0x80002b94
    mem[2790] <= 16'h01d5; // 0x80002b98
    mem[2791] <= 16'h01c7; // 0x80002b9c
    mem[2792] <= 16'hf2e5; // 0x80002ba0
    mem[2793] <= 16'hfff7; // 0x80002ba4
    mem[2794] <= 16'h0000; // 0x80002ba8
    mem[2795] <= 16'hf1df; // 0x80002bac
    mem[2796] <= 16'heb17; // 0x80002bb0
    mem[2797] <= 16'hffee; // 0x80002bb4
    mem[2798] <= 16'h0107; // 0x80002bb8
    mem[2799] <= 16'heb1f; // 0x80002bbc
    mem[2800] <= 16'he6f6; // 0x80002bc0
    mem[2801] <= 16'hffe3; // 0x80002bc4
    mem[2802] <= 16'h0106; // 0x80002bc8
    mem[2803] <= 16'he6df; // 0x80002bcc
    mem[2804] <= 16'h0006; // 0x80002bd0
    mem[2805] <= 16'hf91f; // 0x80002bd4
    mem[2806] <= 16'h0006; // 0x80002bd8
    mem[2807] <= 16'hf4df; // 0x80002bdc
    mem[2808] <= 16'hffe6; // 0x80002be0
    mem[2809] <= 16'h0117; // 0x80002be4
    mem[2810] <= 16'hd6df; // 0x80002be8
    mem[2811] <= 16'hffe7; // 0x80002bec
    mem[2812] <= 16'h0118; // 0x80002bf0
    mem[2813] <= 16'hc31f; // 0x80002bf4
    mem[2814] <= 16'h0006; // 0x80002bf8
    mem[2815] <= 16'h0006; // 0x80002bfc
    mem[2816] <= 16'h0005; // 0x80002c00
    mem[2817] <= 16'h0005; // 0x80002c04
    mem[2818] <= 16'h0c06; // 0x80002c08
    mem[2819] <= 16'h12c5; // 0x80002c0c
    mem[2820] <= 16'h0001; // 0x80002c10
    mem[2821] <= 16'h1ef6; // 0x80002c14
    mem[2822] <= 16'h0100; // 0x80002c18
    mem[2823] <= 16'h0180; // 0x80002c1c
    mem[2824] <= 16'h00f6; // 0x80002c20
    mem[2825] <= 16'h0100; // 0x80002c24
    mem[2826] <= 16'h8000; // 0x80002c28
    mem[2827] <= 16'h0116; // 0x80002c2c
    mem[2828] <= 16'h3407; // 0x80002c30
    mem[2829] <= 16'h00e7; // 0x80002c34
    mem[2830] <= 16'h0007; // 0x80002c38
    mem[2831] <= 16'h0200; // 0x80002c3c
    mem[2832] <= 16'h0117; // 0x80002c40
    mem[2833] <= 16'h411e; // 0x80002c44
    mem[2834] <= 16'h000e; // 0x80002c48
    mem[2835] <= 16'h01c5; // 0x80002c4c
    mem[2836] <= 16'h0115; // 0x80002c50
    mem[2837] <= 16'h01c6; // 0x80002c54
    mem[2838] <= 16'h00b8; // 0x80002c58
    mem[2839] <= 16'h01c5; // 0x80002c5c
    mem[2840] <= 16'h0108; // 0x80002c60
    mem[2841] <= 16'h02c3; // 0x80002c64
    mem[2842] <= 16'h0108; // 0x80002c68
    mem[2843] <= 16'h0105; // 0x80002c6c
    mem[2844] <= 16'h010e; // 0x80002c70
    mem[2845] <= 16'h02c3; // 0x80002c74
    mem[2846] <= 16'h02f5; // 0x80002c78
    mem[2847] <= 16'h0106; // 0x80002c7c
    mem[2848] <= 16'h00e6; // 0x80002c80
    mem[2849] <= 16'h00f7; // 0x80002c84
    mem[2850] <= 16'h0107; // 0x80002c88
    mem[2851] <= 16'h0107; // 0x80002c8c
    mem[2852] <= 16'h36f7; // 0x80002c90
    mem[2853] <= 16'h40f7; // 0x80002c94
    mem[2854] <= 16'h02c7; // 0x80002c98
    mem[2855] <= 16'h010e; // 0x80002c9c
    mem[2856] <= 16'h0107; // 0x80002ca0
    mem[2857] <= 16'h02c7; // 0x80002ca4
    mem[2858] <= 16'h02d5; // 0x80002ca8
    mem[2859] <= 16'h0107; // 0x80002cac
    mem[2860] <= 16'h00f7; // 0x80002cb0
    mem[2861] <= 16'h00a7; // 0x80002cb4
    mem[2862] <= 16'h0107; // 0x80002cb8
    mem[2863] <= 16'h0107; // 0x80002cbc
    mem[2864] <= 16'h00a7; // 0x80002cc0
    mem[2865] <= 16'h0107; // 0x80002cc4
    mem[2866] <= 16'h40a7; // 0x80002cc8
    mem[2867] <= 16'h01c5; // 0x80002ccc
    mem[2868] <= 16'h0000; // 0x80002cd0
    mem[2869] <= 16'h0000; // 0x80002cd4
    mem[2870] <= 16'hfed5; // 0x80002cd8
    mem[2871] <= 16'h0001; // 0x80002cdc
    mem[2872] <= 16'h10f6; // 0x80002ce0
    mem[2873] <= 16'h0100; // 0x80002ce4
    mem[2874] <= 16'h0180; // 0x80002ce8
    mem[2875] <= 16'h00e6; // 0x80002cec
    mem[2876] <= 16'h0100; // 0x80002cf0
    mem[2877] <= 16'h8000; // 0x80002cf4
    mem[2878] <= 16'h340e; // 0x80002cf8
    mem[2879] <= 16'h00f6; // 0x80002cfc
    mem[2880] <= 16'h01c7; // 0x80002d00
    mem[2881] <= 16'h0007; // 0x80002d04
    mem[2882] <= 16'h0200; // 0x80002d08
    mem[2883] <= 16'h00ff; // 0x80002d0c
    mem[2884] <= 16'h41ee; // 0x80002d10
    mem[2885] <= 16'h100e; // 0x80002d14
    mem[2886] <= 16'h0068; // 0x80002d18
    mem[2887] <= 16'h0005; // 0x80002d1c
    mem[2888] <= 16'h010e; // 0x80002d20
    mem[2889] <= 16'h40c5; // 0x80002d24
    mem[2890] <= 16'h40d5; // 0x80002d28
    mem[2891] <= 16'h00f5; // 0x80002d2c
    mem[2892] <= 16'h40d5; // 0x80002d30
    mem[2893] <= 16'h0007; // 0x80002d34
    mem[2894] <= 16'h0003; // 0x80002d38
    mem[2895] <= 16'h0000; // 0x80002d3c
    mem[2896] <= 16'h0006; // 0x80002d40
    mem[2897] <= 16'h0010; // 0x80002d44
    mem[2898] <= 16'h02c8; // 0x80002d48
    mem[2899] <= 16'h0001; // 0x80002d4c
    mem[2900] <= 16'h0af8; // 0x80002d50
    mem[2901] <= 16'h0100; // 0x80002d54
    mem[2902] <= 16'h0180; // 0x80002d58
    mem[2903] <= 16'h00f8; // 0x80002d5c
    mem[2904] <= 16'h0100; // 0x80002d60
    mem[2905] <= 16'h8000; // 0x80002d64
    mem[2906] <= 16'h0118; // 0x80002d68
    mem[2907] <= 16'h3407; // 0x80002d6c
    mem[2908] <= 16'h00e7; // 0x80002d70
    mem[2909] <= 16'h0007; // 0x80002d74
    mem[2910] <= 16'h0200; // 0x80002d78
    mem[2911] <= 16'h0117; // 0x80002d7c
    mem[2912] <= 16'h411e; // 0x80002d80
    mem[2913] <= 16'h1c0e; // 0x80002d84
    mem[2914] <= 16'h0108; // 0x80002d88
    mem[2915] <= 16'h4105; // 0x80002d8c
    mem[2916] <= 16'h0108; // 0x80002d90
    mem[2917] <= 16'h0107; // 0x80002d94
    mem[2918] <= 16'h010e; // 0x80002d98
    mem[2919] <= 16'h02c5; // 0x80002d9c
    mem[2920] <= 16'h02c5; // 0x80002da0
    mem[2921] <= 16'h02f6; // 0x80002da4
    mem[2922] <= 16'h0105; // 0x80002da8
    mem[2923] <= 16'h00e5; // 0x80002dac
    mem[2924] <= 16'h00d7; // 0x80002db0
    mem[2925] <= 16'h0107; // 0x80002db4
    mem[2926] <= 16'h0107; // 0x80002db8
    mem[2927] <= 16'h00d7; // 0x80002dbc
    mem[2928] <= 16'h0107; // 0x80002dc0
    mem[2929] <= 16'h40d7; // 0x80002dc4
    mem[2930] <= 16'h02c7; // 0x80002dc8
    mem[2931] <= 16'h010e; // 0x80002dcc
    mem[2932] <= 16'h010e; // 0x80002dd0
    mem[2933] <= 16'h02c7; // 0x80002dd4
    mem[2934] <= 16'h02f5; // 0x80002dd8
    mem[2935] <= 16'h0107; // 0x80002ddc
    mem[2936] <= 16'h01d7; // 0x80002de0
    mem[2937] <= 16'heea7; // 0x80002de4
    mem[2938] <= 16'hed1f; // 0x80002de8
    mem[2939] <= 16'h0ff0; // 0x80002dec
    mem[2940] <= 16'h00df; // 0x80002df0
    mem[2941] <= 16'h0037; // 0x80002df4
    mem[2942] <= 16'hefdf; // 0x80002df8
    mem[2943] <= 16'h0ff0; // 0x80002dfc
    mem[2944] <= 16'hf707; // 0x80002e00
    mem[2945] <= 16'h0080; // 0x80002e04
    mem[2946] <= 16'hf5df; // 0x80002e08
    mem[2947] <= 16'h0ff0; // 0x80002e0c
    mem[2948] <= 16'he0c7; // 0x80002e10
    mem[2949] <= 16'h0080; // 0x80002e14
    mem[2950] <= 16'he11f; // 0x80002e18
    mem[2951] <= 16'h01e6; // 0x80002e1c
    mem[2952] <= 16'h01c6; // 0x80002e20
    mem[2953] <= 16'h00d7; // 0x80002e24
    mem[2954] <= 16'h01e5; // 0x80002e28
    mem[2955] <= 16'h0106; // 0x80002e2c
    mem[2956] <= 16'h02e8; // 0x80002e30
    mem[2957] <= 16'h0106; // 0x80002e34
    mem[2958] <= 16'h01e5; // 0x80002e38
    mem[2959] <= 16'h010f; // 0x80002e3c
    mem[2960] <= 16'h01c5; // 0x80002e40
    mem[2961] <= 16'h00b7; // 0x80002e44
    mem[2962] <= 16'h01c6; // 0x80002e48
    mem[2963] <= 16'h0105; // 0x80002e4c
    mem[2964] <= 16'h01c5; // 0x80002e50
    mem[2965] <= 16'h02e8; // 0x80002e54
    mem[2966] <= 16'h026f; // 0x80002e58
    mem[2967] <= 16'h0108; // 0x80002e5c
    mem[2968] <= 16'h0108; // 0x80002e60
    mem[2969] <= 16'h00c8; // 0x80002e64
    mem[2970] <= 16'h00d8; // 0x80002e68
    mem[2971] <= 16'hfff3; // 0x80002e6c
    mem[2972] <= 16'h18d8; // 0x80002e70
    mem[2973] <= 16'h0008; // 0x80002e74
    mem[2974] <= 16'h40c8; // 0x80002e78
    mem[2975] <= 16'h02e8; // 0x80002e7c
    mem[2976] <= 16'h0105; // 0x80002e80
    mem[2977] <= 16'h0105; // 0x80002e84
    mem[2978] <= 16'h02e8; // 0x80002e88
    mem[2979] <= 16'h02cf; // 0x80002e8c
    mem[2980] <= 16'h0108; // 0x80002e90
    mem[2981] <= 16'h00b7; // 0x80002e94
    mem[2982] <= 16'h01f7; // 0x80002e98
    mem[2983] <= 16'h00d7; // 0x80002e9c
    mem[2984] <= 16'hfff6; // 0x80002ea0
    mem[2985] <= 16'h14d7; // 0x80002ea4
    mem[2986] <= 16'h0005; // 0x80002ea8
    mem[2987] <= 16'h0103; // 0x80002eac
    mem[2988] <= 16'h0001; // 0x80002eb0
    mem[2989] <= 16'h00c3; // 0x80002eb4
    mem[2990] <= 16'hfff5; // 0x80002eb8
    mem[2991] <= 16'h0113; // 0x80002ebc
    mem[2992] <= 16'h0107; // 0x80002ec0
    mem[2993] <= 16'h0103; // 0x80002ec4
    mem[2994] <= 16'h0117; // 0x80002ec8
    mem[2995] <= 16'h031e; // 0x80002ecc
    mem[2996] <= 16'h41f7; // 0x80002ed0
    mem[2997] <= 16'h02ce; // 0x80002ed4
    mem[2998] <= 16'h0102; // 0x80002ed8
    mem[2999] <= 16'h0313; // 0x80002edc
    mem[3000] <= 16'h011e; // 0x80002ee0
    mem[3001] <= 16'h01d8; // 0x80002ee4
    mem[3002] <= 16'h02c3; // 0x80002ee8
    mem[3003] <= 16'h0118; // 0x80002eec
    mem[3004] <= 16'h00b6; // 0x80002ef0
    mem[3005] <= 16'h0001; // 0x80002ef4
    mem[3006] <= 16'hfff8; // 0x80002ef8
    mem[3007] <= 16'h0108; // 0x80002efc
    mem[3008] <= 16'h0118; // 0x80002f00
    mem[3009] <= 16'h0108; // 0x80002f04
    mem[3010] <= 16'h0112; // 0x80002f08
    mem[3011] <= 16'h00c5; // 0x80002f0c
    mem[3012] <= 16'h0058; // 0x80002f10
    mem[3013] <= 16'h0ac7; // 0x80002f14
    mem[3014] <= 16'h0ec7; // 0x80002f18
    mem[3015] <= 16'h40c7; // 0x80002f1c
    mem[3016] <= 16'h0008; // 0x80002f20
    mem[3017] <= 16'h40f5; // 0x80002f24
    mem[3018] <= 16'h00f5; // 0x80002f28
    mem[3019] <= 16'h40a5; // 0x80002f2c
    mem[3020] <= 16'h01e5; // 0x80002f30
    mem[3021] <= 16'h01c7; // 0x80002f34
    mem[3022] <= 16'h00af; // 0x80002f38
    mem[3023] <= 16'h01c5; // 0x80002f3c
    mem[3024] <= 16'h0000; // 0x80002f40
    mem[3025] <= 16'h01c8; // 0x80002f44
    mem[3026] <= 16'h0115; // 0x80002f48
    mem[3027] <= 16'h0108; // 0x80002f4c
    mem[3028] <= 16'h02c7; // 0x80002f50
    mem[3029] <= 16'h0108; // 0x80002f54
    mem[3030] <= 16'h0107; // 0x80002f58
    mem[3031] <= 16'h0115; // 0x80002f5c
    mem[3032] <= 16'h01c5; // 0x80002f60
    mem[3033] <= 16'h01c5; // 0x80002f64
    mem[3034] <= 16'h00b8; // 0x80002f68
    mem[3035] <= 16'h0105; // 0x80002f6c
    mem[3036] <= 16'h02c7; // 0x80002f70
    mem[3037] <= 16'h02d7; // 0x80002f74
    mem[3038] <= 16'h0107; // 0x80002f78
    mem[3039] <= 16'h0116; // 0x80002f7c
    mem[3040] <= 16'h00a6; // 0x80002f80
    mem[3041] <= 16'h0106; // 0x80002f84
    mem[3042] <= 16'h0106; // 0x80002f88
    mem[3043] <= 16'h00a6; // 0x80002f8c
    mem[3044] <= 16'h0106; // 0x80002f90
    mem[3045] <= 16'h40a6; // 0x80002f94
    mem[3046] <= 16'h02c6; // 0x80002f98
    mem[3047] <= 16'h0105; // 0x80002f9c
    mem[3048] <= 16'h0108; // 0x80002fa0
    mem[3049] <= 16'h02c6; // 0x80002fa4
    mem[3050] <= 16'h02e7; // 0x80002fa8
    mem[3051] <= 16'h0106; // 0x80002fac
    mem[3052] <= 16'h0115; // 0x80002fb0
    mem[3053] <= 16'h00e5; // 0x80002fb4
    mem[3054] <= 16'h0105; // 0x80002fb8
    mem[3055] <= 16'h0105; // 0x80002fbc
    mem[3056] <= 16'h00e5; // 0x80002fc0
    mem[3057] <= 16'h0105; // 0x80002fc4
    mem[3058] <= 16'h40e5; // 0x80002fc8
    mem[3059] <= 16'hdcdf; // 0x80002fcc
    mem[3060] <= 16'h40f8; // 0x80002fd0
    mem[3061] <= 16'h40d6; // 0x80002fd4
    mem[3062] <= 16'h00f8; // 0x80002fd8
    mem[3063] <= 16'h4105; // 0x80002fdc
    mem[3064] <= 16'h40b7; // 0x80002fe0
    mem[3065] <= 16'hf41f; // 0x80002fe4
    mem[3066] <= 16'hedf7; // 0x80002fe8
    mem[3067] <= 16'hffe6; // 0x80002fec
    mem[3068] <= 16'h00d7; // 0x80002ff0
    mem[3069] <= 16'heb9f; // 0x80002ff4
    mem[3070] <= 16'he6c8; // 0x80002ff8
    mem[3071] <= 16'hffe3; // 0x80002ffc
    mem[3072] <= 16'h00d8; // 0x80003000
    mem[3073] <= 16'he75f; // 0x80003004
    mem[3074] <= 16'h0107; // 0x80003008
    mem[3075] <= 16'hc89f; // 0x8000300c
    mem[3076] <= 16'hfd05; // 0x80003010
    mem[3077] <= 16'h0008; // 0x80003014
    mem[3078] <= 16'h0000; // 0x80003018
    mem[3079] <= 16'hf09f; // 0x8000301c
    mem[3080] <= 16'h0005; // 0x80003020
    mem[3081] <= 16'h0000; // 0x80003024
    mem[3082] <= 16'h0015; // 0x80003028
    mem[3083] <= 16'h0006; // 0x8000302c
    mem[3084] <= 16'h00c5; // 0x80003030
    mem[3085] <= 16'h0015; // 0x80003034
    mem[3086] <= 16'h0016; // 0x80003038
    mem[3087] <= 16'hfe05; // 0x8000303c
    mem[3088] <= 16'h0000; // 0x80003040
 
 
//================================================================
//== Section  .text.startup
//================================================================
    mem[3089] <= 16'h2000; // 0x80003044
    mem[3090] <= 16'h0020; // 0x80003048
    mem[3091] <= 16'h0007; // 0x8000304c
    mem[3092] <= 16'hfed7; // 0x80003050
    mem[3093] <= 16'h0040; // 0x80003054
    mem[3094] <= 16'h00e7; // 0x80003058
    mem[3095] <= 16'h0800; // 0x8000305c
    mem[3096] <= 16'h3047; // 0x80003060
    mem[3097] <= 16'h0000; // 0x80003064
    mem[3098] <= 16'hff01; // 0x80003068
    mem[3099] <= 16'h0000; // 0x8000306c
    mem[3100] <= 16'h3e85; // 0x80003070
    mem[3101] <= 16'h0011; // 0x80003074
    mem[3102] <= 16'hffff; // 0x80003078
    mem[3103] <= 16'ha4c3; // 0x8000307c
    mem[3104] <= 16'h00c1; // 0x80003080
    mem[3105] <= 16'hfff0; // 0x80003084
    mem[3106] <= 16'h0101; // 0x80003088
    mem[3107] <= 16'h0000; // 0x8000308c
 
 
//================================================================
//== Section  .rodata
//================================================================
    mem[3108] <= 16'hffff; // 0x80003090
    mem[3109] <= 16'hffff; // 0x80003094
    mem[3110] <= 16'hffff; // 0x80003098
    mem[3111] <= 16'hffff; // 0x8000309c
    mem[3112] <= 16'hffff; // 0x800030a0
    mem[3113] <= 16'hffff; // 0x800030a4
    mem[3114] <= 16'hffff; // 0x800030a8
    mem[3115] <= 16'hffff; // 0x800030ac
    mem[3116] <= 16'hffff; // 0x800030b0
    mem[3117] <= 16'hffff; // 0x800030b4
    mem[3118] <= 16'hffff; // 0x800030b8
    mem[3119] <= 16'hffff; // 0x800030bc
    mem[3120] <= 16'hffff; // 0x800030c0
    mem[3121] <= 16'hffff; // 0x800030c4
    mem[3122] <= 16'hffff; // 0x800030c8
    mem[3123] <= 16'hffff; // 0x800030cc
    mem[3124] <= 16'hffff; // 0x800030d0
    mem[3125] <= 16'hffff; // 0x800030d4
    mem[3126] <= 16'hffff; // 0x800030d8
    mem[3127] <= 16'hffff; // 0x800030dc
    mem[3128] <= 16'hffff; // 0x800030e0
    mem[3129] <= 16'hffff; // 0x800030e4
    mem[3130] <= 16'hffff; // 0x800030e8
    mem[3131] <= 16'hffff; // 0x800030ec
    mem[3132] <= 16'hffff; // 0x800030f0
    mem[3133] <= 16'hffff; // 0x800030f4
    mem[3134] <= 16'hffff; // 0x800030f8
    mem[3135] <= 16'hffff; // 0x800030fc
    mem[3136] <= 16'hffff; // 0x80003100
    mem[3137] <= 16'hffff; // 0x80003104
    mem[3138] <= 16'hffff; // 0x80003108
    mem[3139] <= 16'hffff; // 0x8000310c
    mem[3140] <= 16'hffff; // 0x80003110
    mem[3141] <= 16'hffff; // 0x80003114
    mem[3142] <= 16'hffff; // 0x80003118
    mem[3143] <= 16'hffff; // 0x8000311c
    mem[3144] <= 16'hffff; // 0x80003120
    mem[3145] <= 16'hffff; // 0x80003124
    mem[3146] <= 16'hffff; // 0x80003128
    mem[3147] <= 16'hffff; // 0x8000312c
    mem[3148] <= 16'hffff; // 0x80003130
    mem[3149] <= 16'hffff; // 0x80003134
    mem[3150] <= 16'hffff; // 0x80003138
    mem[3151] <= 16'hffff; // 0x8000313c
    mem[3152] <= 16'hffff; // 0x80003140
    mem[3153] <= 16'hffff; // 0x80003144
    mem[3154] <= 16'hffff; // 0x80003148
    mem[3155] <= 16'hffff; // 0x8000314c
    mem[3156] <= 16'hffff; // 0x80003150
    mem[3157] <= 16'hffff; // 0x80003154
    mem[3158] <= 16'hffff; // 0x80003158
    mem[3159] <= 16'hffff; // 0x8000315c
    mem[3160] <= 16'hffff; // 0x80003160
    mem[3161] <= 16'hffff; // 0x80003164
    mem[3162] <= 16'hffff; // 0x80003168
    mem[3163] <= 16'hffff; // 0x8000316c
    mem[3164] <= 16'hffff; // 0x80003170
    mem[3165] <= 16'hffff; // 0x80003174
    mem[3166] <= 16'hffff; // 0x80003178
    mem[3167] <= 16'hffff; // 0x8000317c
    mem[3168] <= 16'hffff; // 0x80003180
    mem[3169] <= 16'hffff; // 0x80003184
    mem[3170] <= 16'hffff; // 0x80003188
    mem[3171] <= 16'hffff; // 0x8000318c
    mem[3172] <= 16'hffff; // 0x80003190
    mem[3173] <= 16'hffff; // 0x80003194
    mem[3174] <= 16'hffff; // 0x80003198
    mem[3175] <= 16'hffff; // 0x8000319c
    mem[3176] <= 16'hffff; // 0x800031a0
    mem[3177] <= 16'hffff; // 0x800031a4
    mem[3178] <= 16'hffff; // 0x800031a8
    mem[3179] <= 16'hffff; // 0x800031ac
    mem[3180] <= 16'hffff; // 0x800031b0
    mem[3181] <= 16'hffff; // 0x800031b4
    mem[3182] <= 16'hffff; // 0x800031b8
    mem[3183] <= 16'hffff; // 0x800031bc
    mem[3184] <= 16'hffff; // 0x800031c0
    mem[3185] <= 16'hffff; // 0x800031c4
    mem[3186] <= 16'hffff; // 0x800031c8
    mem[3187] <= 16'hffff; // 0x800031cc
    mem[3188] <= 16'hffff; // 0x800031d0
    mem[3189] <= 16'hffff; // 0x800031d4
    mem[3190] <= 16'hffff; // 0x800031d8
    mem[3191] <= 16'hffff; // 0x800031dc
    mem[3192] <= 16'hffff; // 0x800031e0
    mem[3193] <= 16'hffff; // 0x800031e4
    mem[3194] <= 16'hffff; // 0x800031e8
    mem[3195] <= 16'hffff; // 0x800031ec
    mem[3196] <= 16'hffff; // 0x800031f0
    mem[3197] <= 16'hffff; // 0x800031f4
    mem[3198] <= 16'hffff; // 0x800031f8
    mem[3199] <= 16'hffff; // 0x800031fc
    mem[3200] <= 16'hffff; // 0x80003200
    mem[3201] <= 16'hffff; // 0x80003204
    mem[3202] <= 16'hffff; // 0x80003208
    mem[3203] <= 16'hffff; // 0x8000320c
    mem[3204] <= 16'hffff; // 0x80003210
    mem[3205] <= 16'hffff; // 0x80003214
    mem[3206] <= 16'hffff; // 0x80003218
    mem[3207] <= 16'hffff; // 0x8000321c
    mem[3208] <= 16'hffff; // 0x80003220
    mem[3209] <= 16'hffff; // 0x80003224
    mem[3210] <= 16'hffff; // 0x80003228
    mem[3211] <= 16'hffff; // 0x8000322c
    mem[3212] <= 16'hffff; // 0x80003230
    mem[3213] <= 16'hffff; // 0x80003234
    mem[3214] <= 16'hffff; // 0x80003238
    mem[3215] <= 16'hffff; // 0x8000323c
    mem[3216] <= 16'hffff; // 0x80003240
    mem[3217] <= 16'hffff; // 0x80003244
    mem[3218] <= 16'hffff; // 0x80003248
    mem[3219] <= 16'hffff; // 0x8000324c
    mem[3220] <= 16'hffff; // 0x80003250
    mem[3221] <= 16'hffff; // 0x80003254
    mem[3222] <= 16'hffff; // 0x80003258
    mem[3223] <= 16'hffff; // 0x8000325c
    mem[3224] <= 16'hffff; // 0x80003260
    mem[3225] <= 16'hffff; // 0x80003264
    mem[3226] <= 16'hffff; // 0x80003268
    mem[3227] <= 16'hffff; // 0x8000326c
    mem[3228] <= 16'hffff; // 0x80003270
    mem[3229] <= 16'hffff; // 0x80003274
    mem[3230] <= 16'hffff; // 0x80003278
    mem[3231] <= 16'hffff; // 0x8000327c
    mem[3232] <= 16'hffff; // 0x80003280
    mem[3233] <= 16'hffff; // 0x80003284
    mem[3234] <= 16'hffff; // 0x80003288
    mem[3235] <= 16'hffff; // 0x8000328c
    mem[3236] <= 16'hffff; // 0x80003290
    mem[3237] <= 16'hffff; // 0x80003294
    mem[3238] <= 16'hffff; // 0x80003298
    mem[3239] <= 16'hffff; // 0x8000329c
    mem[3240] <= 16'hffff; // 0x800032a0
    mem[3241] <= 16'hffff; // 0x800032a4
    mem[3242] <= 16'hffff; // 0x800032a8
    mem[3243] <= 16'hffff; // 0x800032ac
    mem[3244] <= 16'hffff; // 0x800032b0
    mem[3245] <= 16'hffff; // 0x800032b4
    mem[3246] <= 16'hffff; // 0x800032b8
    mem[3247] <= 16'hffff; // 0x800032bc
    mem[3248] <= 16'hffff; // 0x800032c0
    mem[3249] <= 16'hffff; // 0x800032c4
    mem[3250] <= 16'hffff; // 0x800032c8
    mem[3251] <= 16'hffff; // 0x800032cc
    mem[3252] <= 16'hffff; // 0x800032d0
    mem[3253] <= 16'hffff; // 0x800032d4
    mem[3254] <= 16'hffff; // 0x800032d8
    mem[3255] <= 16'hffff; // 0x800032dc
    mem[3256] <= 16'hffff; // 0x800032e0
    mem[3257] <= 16'hffff; // 0x800032e4
    mem[3258] <= 16'hffff; // 0x800032e8
    mem[3259] <= 16'hffff; // 0x800032ec
    mem[3260] <= 16'hffff; // 0x800032f0
    mem[3261] <= 16'hffff; // 0x800032f4
    mem[3262] <= 16'hffff; // 0x800032f8
    mem[3263] <= 16'hffff; // 0x800032fc
    mem[3264] <= 16'hffff; // 0x80003300
    mem[3265] <= 16'hffff; // 0x80003304
    mem[3266] <= 16'hffff; // 0x80003308
    mem[3267] <= 16'hffff; // 0x8000330c
    mem[3268] <= 16'hffff; // 0x80003310
    mem[3269] <= 16'hffff; // 0x80003314
    mem[3270] <= 16'hffff; // 0x80003318
    mem[3271] <= 16'hffff; // 0x8000331c
    mem[3272] <= 16'hffff; // 0x80003320
    mem[3273] <= 16'hffff; // 0x80003324
    mem[3274] <= 16'hffff; // 0x80003328
    mem[3275] <= 16'hffff; // 0x8000332c
    mem[3276] <= 16'hffff; // 0x80003330
    mem[3277] <= 16'hffff; // 0x80003334
    mem[3278] <= 16'hffff; // 0x80003338
    mem[3279] <= 16'hffff; // 0x8000333c
    mem[3280] <= 16'h0202; // 0x80003340
    mem[3281] <= 16'h0303; // 0x80003344
    mem[3282] <= 16'h0404; // 0x80003348
    mem[3283] <= 16'h0404; // 0x8000334c
    mem[3284] <= 16'h0505; // 0x80003350
    mem[3285] <= 16'h0505; // 0x80003354
    mem[3286] <= 16'h0505; // 0x80003358
    mem[3287] <= 16'h0505; // 0x8000335c
    mem[3288] <= 16'h0606; // 0x80003360
    mem[3289] <= 16'h0606; // 0x80003364
    mem[3290] <= 16'h0606; // 0x80003368
    mem[3291] <= 16'h0606; // 0x8000336c
    mem[3292] <= 16'h0606; // 0x80003370
    mem[3293] <= 16'h0606; // 0x80003374
    mem[3294] <= 16'h0606; // 0x80003378
    mem[3295] <= 16'h0606; // 0x8000337c
    mem[3296] <= 16'h0707; // 0x80003380
    mem[3297] <= 16'h0707; // 0x80003384
    mem[3298] <= 16'h0707; // 0x80003388
    mem[3299] <= 16'h0707; // 0x8000338c
    mem[3300] <= 16'h0707; // 0x80003390
    mem[3301] <= 16'h0707; // 0x80003394
    mem[3302] <= 16'h0707; // 0x80003398
    mem[3303] <= 16'h0707; // 0x8000339c
    mem[3304] <= 16'h0707; // 0x800033a0
    mem[3305] <= 16'h0707; // 0x800033a4
    mem[3306] <= 16'h0707; // 0x800033a8
    mem[3307] <= 16'h0707; // 0x800033ac
    mem[3308] <= 16'h0707; // 0x800033b0
    mem[3309] <= 16'h0707; // 0x800033b4
    mem[3310] <= 16'h0707; // 0x800033b8
    mem[3311] <= 16'h0707; // 0x800033bc
    mem[3312] <= 16'h0808; // 0x800033c0
    mem[3313] <= 16'h0808; // 0x800033c4
    mem[3314] <= 16'h0808; // 0x800033c8
    mem[3315] <= 16'h0808; // 0x800033cc
    mem[3316] <= 16'h0808; // 0x800033d0
    mem[3317] <= 16'h0808; // 0x800033d4
    mem[3318] <= 16'h0808; // 0x800033d8
    mem[3319] <= 16'h0808; // 0x800033dc
    mem[3320] <= 16'h0808; // 0x800033e0
    mem[3321] <= 16'h0808; // 0x800033e4
    mem[3322] <= 16'h0808; // 0x800033e8
    mem[3323] <= 16'h0808; // 0x800033ec
    mem[3324] <= 16'h0808; // 0x800033f0
    mem[3325] <= 16'h0808; // 0x800033f4
    mem[3326] <= 16'h0808; // 0x800033f8
    mem[3327] <= 16'h0808; // 0x800033fc
    mem[3328] <= 16'h0808; // 0x80003400
    mem[3329] <= 16'h0808; // 0x80003404
    mem[3330] <= 16'h0808; // 0x80003408
    mem[3331] <= 16'h0808; // 0x8000340c
    mem[3332] <= 16'h0808; // 0x80003410
    mem[3333] <= 16'h0808; // 0x80003414
    mem[3334] <= 16'h0808; // 0x80003418
    mem[3335] <= 16'h0808; // 0x8000341c
    mem[3336] <= 16'h0808; // 0x80003420
    mem[3337] <= 16'h0808; // 0x80003424
    mem[3338] <= 16'h0808; // 0x80003428
    mem[3339] <= 16'h0808; // 0x8000342c
    mem[3340] <= 16'h0808; // 0x80003430
    mem[3341] <= 16'h0808; // 0x80003434
    mem[3342] <= 16'h0808; // 0x80003438
    mem[3343] <= 16'h0808; // 0x8000343c
 
 
//================================================================
//== Section  .rodata.str1.4
//================================================================
    mem[3344] <= 16'h6379; // 0x80003440
    mem[3345] <= 16'h0000; // 0x80003444
    mem[3346] <= 16'h736e; // 0x80003448
    mem[3347] <= 16'h7465; // 0x8000344c
    mem[3348] <= 16'h0000; // 0x80003450
    mem[3349] <= 16'h6c70; // 0x80003454
    mem[3350] <= 16'h6e65; // 0x80003458
    mem[3351] <= 16'h616d; // 0x8000345c
    mem[3352] <= 16'h2928; // 0x80003460
    mem[3353] <= 16'h6f66; // 0x80003464
    mem[3354] <= 16'h000a; // 0x80003468
    mem[3355] <= 16'h6c75; // 0x8000346c
    mem[3356] <= 16'h0000; // 0x80003470
    mem[3357] <= 16'h3d20; // 0x80003474
    mem[3358] <= 16'h0a64; // 0x80003478
    mem[3359] <= 16'h0000; // 0x8000347c
 
 
//================================================================
//== Section  .eh_frame
//================================================================
    mem[3360] <= 16'h0000; // 0x80003480
    mem[3361] <= 16'h0000; // 0x80003484
    mem[3362] <= 16'h0052; // 0x80003488
    mem[3363] <= 16'h0101; // 0x8000348c
    mem[3364] <= 16'h0002; // 0x80003490
    mem[3365] <= 16'h0000; // 0x80003494
    mem[3366] <= 16'h0000; // 0x80003498
    mem[3367] <= 16'hffff; // 0x8000349c
    mem[3368] <= 16'h0000; // 0x800034a0
    mem[3369] <= 16'h0000; // 0x800034a4
    mem[3370] <= 16'h0000; // 0x800034a8
    mem[3371] <= 16'h0000; // 0x800034ac
    mem[3372] <= 16'hffff; // 0x800034b0
    mem[3373] <= 16'h0000; // 0x800034b4
    mem[3374] <= 16'h0000; // 0x800034b8
 
 
end
endmodule
 
 
 
module single_port_ram_sim_low #(parameter ADDR_WIDTH, DATA_WIDTH ) (
    input  wire [ADDR_WIDTH - 1 : 0]         addr,
    input  wire [DATA_WIDTH - 1 : 0]         din,
    input  wire [DATA_WIDTH / 8 - 1 : 0]     write_en,
    input  wire                              clk,
    output reg [DATA_WIDTH - 1 : 0]          dout
);
    reg [DATA_WIDTH - 1 : 0] mem [(1<<ADDR_WIDTH)-1:0];
    genvar i;
    generate
        for (i = 0; i < (DATA_WIDTH / 8); i = i + 1) begin : gen_proc
            always @(posedge clk) begin
                if (write_en[i]) begin
                    mem[(addr)][8 * (i + 1) - 1 : 8 * i] <= din[8 * (i + 1) - 1 : 8 * i];
                end
            end
        end
    endgenerate
 
    always @(posedge clk) begin
        dout <= mem[addr];
    end
 
initial begin
//================================================================
//== Section  .note.gnu.build-id
//================================================================
    mem[0] <= 16'h0004; // 0x80000000
    mem[1] <= 16'h0014; // 0x80000004
    mem[2] <= 16'h0003; // 0x80000008
    mem[3] <= 16'h4e47; // 0x8000000c
    mem[4] <= 16'hf6c7; // 0x80000010
    mem[5] <= 16'hdd30; // 0x80000014
    mem[6] <= 16'h1240; // 0x80000018
    mem[7] <= 16'h3f36; // 0x8000001c
    mem[8] <= 16'h0789; // 0x80000020
 
 
//================================================================
//== Section  .text.init
//================================================================
    mem[9] <= 16'h0093; // 0x80000024
    mem[10] <= 16'h0113; // 0x80000028
    mem[11] <= 16'h0193; // 0x8000002c
    mem[12] <= 16'h0213; // 0x80000030
    mem[13] <= 16'h0293; // 0x80000034
    mem[14] <= 16'h0313; // 0x80000038
    mem[15] <= 16'h0393; // 0x8000003c
    mem[16] <= 16'h0413; // 0x80000040
    mem[17] <= 16'h0493; // 0x80000044
    mem[18] <= 16'h0513; // 0x80000048
    mem[19] <= 16'h0593; // 0x8000004c
    mem[20] <= 16'h0613; // 0x80000050
    mem[21] <= 16'h0693; // 0x80000054
    mem[22] <= 16'h0713; // 0x80000058
    mem[23] <= 16'h0793; // 0x8000005c
    mem[24] <= 16'h0813; // 0x80000060
    mem[25] <= 16'h0893; // 0x80000064
    mem[26] <= 16'h0913; // 0x80000068
    mem[27] <= 16'h0993; // 0x8000006c
    mem[28] <= 16'h0a13; // 0x80000070
    mem[29] <= 16'h0a93; // 0x80000074
    mem[30] <= 16'h0b13; // 0x80000078
    mem[31] <= 16'h0b93; // 0x8000007c
    mem[32] <= 16'h0c13; // 0x80000080
    mem[33] <= 16'h0c93; // 0x80000084
    mem[34] <= 16'h0d13; // 0x80000088
    mem[35] <= 16'h0d93; // 0x8000008c
    mem[36] <= 16'h0e13; // 0x80000090
    mem[37] <= 16'h0e93; // 0x80000094
    mem[38] <= 16'h0f13; // 0x80000098
    mem[39] <= 16'h0f93; // 0x8000009c
    mem[40] <= 16'he2b7; // 0x800000a0
    mem[41] <= 16'ha073; // 0x800000a4
    mem[42] <= 16'h0293; // 0x800000a8
    mem[43] <= 16'h9293; // 0x800000ac
    mem[44] <= 16'hca63; // 0x800000b0
    mem[45] <= 16'h0513; // 0x800000b4
    mem[46] <= 16'h1297; // 0x800000b8
    mem[47] <= 16'ha423; // 0x800000bc
    mem[48] <= 16'hf06f; // 0x800000c0
    mem[49] <= 16'h0297; // 0x800000c4
    mem[50] <= 16'h8293; // 0x800000c8
    mem[51] <= 16'h9073; // 0x800000cc
    mem[52] <= 16'h4197; // 0x800000d0
    mem[53] <= 16'h8193; // 0x800000d4
    mem[54] <= 16'h6217; // 0x800000d8
    mem[55] <= 16'h0213; // 0x800000dc
    mem[56] <= 16'h7213; // 0x800000e0
    mem[57] <= 16'h2573; // 0x800000e4
    mem[58] <= 16'h0593; // 0x800000e8
    mem[59] <= 16'h7063; // 0x800000ec
    mem[60] <= 16'h1613; // 0x800000f0
    mem[61] <= 16'h0233; // 0x800000f4
    mem[62] <= 16'h0113; // 0x800000f8
    mem[63] <= 16'h1113; // 0x800000fc
    mem[64] <= 16'h0133; // 0x80000100
    mem[65] <= 16'h206f; // 0x80000104
    mem[66] <= 16'h0113; // 0x80000108
    mem[67] <= 16'h2223; // 0x8000010c
    mem[68] <= 16'h2423; // 0x80000110
    mem[69] <= 16'h2623; // 0x80000114
    mem[70] <= 16'h2823; // 0x80000118
    mem[71] <= 16'h2a23; // 0x8000011c
    mem[72] <= 16'h2c23; // 0x80000120
    mem[73] <= 16'h2e23; // 0x80000124
    mem[74] <= 16'h2023; // 0x80000128
    mem[75] <= 16'h2223; // 0x8000012c
    mem[76] <= 16'h2423; // 0x80000130
    mem[77] <= 16'h2623; // 0x80000134
    mem[78] <= 16'h2823; // 0x80000138
    mem[79] <= 16'h2a23; // 0x8000013c
    mem[80] <= 16'h2c23; // 0x80000140
    mem[81] <= 16'h2e23; // 0x80000144
    mem[82] <= 16'h2023; // 0x80000148
    mem[83] <= 16'h2223; // 0x8000014c
    mem[84] <= 16'h2423; // 0x80000150
    mem[85] <= 16'h2623; // 0x80000154
    mem[86] <= 16'h2823; // 0x80000158
    mem[87] <= 16'h2a23; // 0x8000015c
    mem[88] <= 16'h2c23; // 0x80000160
    mem[89] <= 16'h2e23; // 0x80000164
    mem[90] <= 16'h2023; // 0x80000168
    mem[91] <= 16'h2223; // 0x8000016c
    mem[92] <= 16'h2423; // 0x80000170
    mem[93] <= 16'h2623; // 0x80000174
    mem[94] <= 16'h2823; // 0x80000178
    mem[95] <= 16'h2a23; // 0x8000017c
    mem[96] <= 16'h2c23; // 0x80000180
    mem[97] <= 16'h2e23; // 0x80000184
    mem[98] <= 16'h2573; // 0x80000188
    mem[99] <= 16'h25f3; // 0x8000018c
    mem[100] <= 16'h0613; // 0x80000190
    mem[101] <= 16'h10ef; // 0x80000194
    mem[102] <= 16'h1073; // 0x80000198
    mem[103] <= 16'h22b7; // 0x8000019c
    mem[104] <= 16'h8293; // 0x800001a0
    mem[105] <= 16'ha073; // 0x800001a4
    mem[106] <= 16'h2083; // 0x800001a8
    mem[107] <= 16'h2103; // 0x800001ac
    mem[108] <= 16'h2183; // 0x800001b0
    mem[109] <= 16'h2203; // 0x800001b4
    mem[110] <= 16'h2283; // 0x800001b8
    mem[111] <= 16'h2303; // 0x800001bc
    mem[112] <= 16'h2383; // 0x800001c0
    mem[113] <= 16'h2403; // 0x800001c4
    mem[114] <= 16'h2483; // 0x800001c8
    mem[115] <= 16'h2503; // 0x800001cc
    mem[116] <= 16'h2583; // 0x800001d0
    mem[117] <= 16'h2603; // 0x800001d4
    mem[118] <= 16'h2683; // 0x800001d8
    mem[119] <= 16'h2703; // 0x800001dc
    mem[120] <= 16'h2783; // 0x800001e0
    mem[121] <= 16'h2803; // 0x800001e4
    mem[122] <= 16'h2883; // 0x800001e8
    mem[123] <= 16'h2903; // 0x800001ec
    mem[124] <= 16'h2983; // 0x800001f0
    mem[125] <= 16'h2a03; // 0x800001f4
    mem[126] <= 16'h2a83; // 0x800001f8
    mem[127] <= 16'h2b03; // 0x800001fc
    mem[128] <= 16'h2b83; // 0x80000200
    mem[129] <= 16'h2c03; // 0x80000204
    mem[130] <= 16'h2c83; // 0x80000208
    mem[131] <= 16'h2d03; // 0x8000020c
    mem[132] <= 16'h2d83; // 0x80000210
    mem[133] <= 16'h2e03; // 0x80000214
    mem[134] <= 16'h2e83; // 0x80000218
    mem[135] <= 16'h2f03; // 0x8000021c
    mem[136] <= 16'h2f83; // 0x80000220
    mem[137] <= 16'h0113; // 0x80000224
    mem[138] <= 16'h0073; // 0x80000228
 
 
//================================================================
//== Section  .tohost
//================================================================
    mem[1024] <= 16'h0000; // 0x80001000
    mem[1025] <= 16'h0000; // 0x80001004
    mem[1026] <= 16'h0000; // 0x80001008
    mem[1027] <= 16'h0000; // 0x8000100c
    mem[1028] <= 16'h0000; // 0x80001010
    mem[1029] <= 16'h0000; // 0x80001014
    mem[1030] <= 16'h0000; // 0x80001018
    mem[1031] <= 16'h0000; // 0x8000101c
    mem[1032] <= 16'h0000; // 0x80001020
    mem[1033] <= 16'h0000; // 0x80001024
    mem[1034] <= 16'h0000; // 0x80001028
    mem[1035] <= 16'h0000; // 0x8000102c
    mem[1036] <= 16'h0000; // 0x80001030
    mem[1037] <= 16'h0000; // 0x80001034
    mem[1038] <= 16'h0000; // 0x80001038
    mem[1039] <= 16'h0000; // 0x8000103c
    mem[1040] <= 16'h0000; // 0x80001040
    mem[1041] <= 16'h0000; // 0x80001044
 
 
//================================================================
//== Section  .text
//================================================================
    mem[1042] <= 16'h0513; // 0x80001048
    mem[1043] <= 16'h05b3; // 0x8000104c
    mem[1044] <= 16'h2023; // 0x80001050
    mem[1045] <= 16'h8067; // 0x80001054
    mem[1046] <= 16'h0113; // 0x80001058
    mem[1047] <= 16'h2623; // 0x8000105c
    mem[1048] <= 16'h0993; // 0x80001060
    mem[1049] <= 16'h2a23; // 0x80001064
    mem[1050] <= 16'h9493; // 0x80001068
    mem[1051] <= 16'h2e23; // 0x8000106c
    mem[1052] <= 16'h2c23; // 0x80001070
    mem[1053] <= 16'h2823; // 0x80001074
    mem[1054] <= 16'h04b3; // 0x80001078
    mem[1055] <= 16'h8413; // 0x8000107c
    mem[1056] <= 16'hac23; // 0x80001080
    mem[1057] <= 16'h0913; // 0x80001084
    mem[1058] <= 16'ha023; // 0x80001088
    mem[1059] <= 16'ha223; // 0x8000108c
    mem[1060] <= 16'h8513; // 0x80001090
    mem[1061] <= 16'h0593; // 0x80001094
    mem[1062] <= 16'h10ef; // 0x80001098
    mem[1063] <= 16'h1913; // 0x8000109c
    mem[1064] <= 16'h07b3; // 0x800010a0
    mem[1065] <= 16'h07b3; // 0x800010a4
    mem[1066] <= 16'ha703; // 0x800010a8
    mem[1067] <= 16'haa23; // 0x800010ac
    mem[1068] <= 16'hac23; // 0x800010b0
    mem[1069] <= 16'h0713; // 0x800010b4
    mem[1070] <= 16'ha823; // 0x800010b8
    mem[1071] <= 16'ha703; // 0x800010bc
    mem[1072] <= 16'h0433; // 0x800010c0
    mem[1073] <= 16'h2083; // 0x800010c4
    mem[1074] <= 16'h0433; // 0x800010c8
    mem[1075] <= 16'h17b7; // 0x800010cc
    mem[1076] <= 16'h8433; // 0x800010d0
    mem[1077] <= 16'h0793; // 0x800010d4
    mem[1078] <= 16'h2a23; // 0x800010d8
    mem[1079] <= 16'h2483; // 0x800010dc
    mem[1080] <= 16'h2403; // 0x800010e0
    mem[1081] <= 16'h2903; // 0x800010e4
    mem[1082] <= 16'h2983; // 0x800010e8
    mem[1083] <= 16'h2297; // 0x800010ec
    mem[1084] <= 16'ha023; // 0x800010f0
    mem[1085] <= 16'h0113; // 0x800010f4
    mem[1086] <= 16'h8067; // 0x800010f8
    mem[1087] <= 16'h7513; // 0x800010fc
    mem[1088] <= 16'hf593; // 0x80001100
    mem[1089] <= 16'h0663; // 0x80001104
    mem[1090] <= 16'h0513; // 0x80001108
    mem[1091] <= 16'h8067; // 0x8000110c
    mem[1092] <= 16'h2297; // 0x80001110
    mem[1093] <= 16'h8aa3; // 0x80001114
    mem[1094] <= 16'h0513; // 0x80001118
    mem[1095] <= 16'h8067; // 0x8000111c
    mem[1096] <= 16'h0113; // 0x80001120
    mem[1097] <= 16'h2423; // 0x80001124
    mem[1098] <= 16'h2223; // 0x80001128
    mem[1099] <= 16'h2623; // 0x8000112c
    mem[1100] <= 16'h0413; // 0x80001130
    mem[1101] <= 16'h8493; // 0x80001134
    mem[1102] <= 16'hc583; // 0x80001138
    mem[1103] <= 16'h4503; // 0x8000113c
    mem[1104] <= 16'hf0ef; // 0x80001140
    mem[1105] <= 16'h1ae3; // 0x80001144
    mem[1106] <= 16'h8593; // 0x80001148
    mem[1107] <= 16'h0513; // 0x8000114c
    mem[1108] <= 16'h10ef; // 0x80001150
    mem[1109] <= 16'h5463; // 0x80001154
    mem[1110] <= 16'h2083; // 0x80001158
    mem[1111] <= 16'h0793; // 0x8000115c
    mem[1112] <= 16'h0513; // 0x80001160
    mem[1113] <= 16'h2403; // 0x80001164
    mem[1114] <= 16'h2483; // 0x80001168
    mem[1115] <= 16'h2297; // 0x8000116c
    mem[1116] <= 16'ha023; // 0x80001170
    mem[1117] <= 16'h0113; // 0x80001174
    mem[1118] <= 16'h8067; // 0x80001178
    mem[1119] <= 16'h2083; // 0x8000117c
    mem[1120] <= 16'h0513; // 0x80001180
    mem[1121] <= 16'h2403; // 0x80001184
    mem[1122] <= 16'h2483; // 0x80001188
    mem[1123] <= 16'h0113; // 0x8000118c
    mem[1124] <= 16'h8067; // 0x80001190
    mem[1125] <= 16'h0513; // 0x80001194
    mem[1126] <= 16'h3513; // 0x80001198
    mem[1127] <= 16'h8067; // 0x8000119c
    mem[1128] <= 16'h0113; // 0x800011a0
    mem[1129] <= 16'h2423; // 0x800011a4
    mem[1130] <= 16'h2223; // 0x800011a8
    mem[1131] <= 16'h2623; // 0x800011ac
    mem[1132] <= 16'h0413; // 0x800011b0
    mem[1133] <= 16'h8493; // 0x800011b4
    mem[1134] <= 16'hf0ef; // 0x800011b8
    mem[1135] <= 16'h0e63; // 0x800011bc
    mem[1136] <= 16'ha023; // 0x800011c0
    mem[1137] <= 16'h0793; // 0x800011c4
    mem[1138] <= 16'h0063; // 0x800011c8
    mem[1139] <= 16'h0663; // 0x800011cc
    mem[1140] <= 16'h0713; // 0x800011d0
    mem[1141] <= 16'h0e63; // 0x800011d4
    mem[1142] <= 16'h0793; // 0x800011d8
    mem[1143] <= 16'h1463; // 0x800011dc
    mem[1144] <= 16'ha023; // 0x800011e0
    mem[1145] <= 16'h2083; // 0x800011e4
    mem[1146] <= 16'h2403; // 0x800011e8
    mem[1147] <= 16'h2483; // 0x800011ec
    mem[1148] <= 16'h0113; // 0x800011f0
    mem[1149] <= 16'h8067; // 0x800011f4
    mem[1150] <= 16'h0793; // 0x800011f8
    mem[1151] <= 16'ha023; // 0x800011fc
    mem[1152] <= 16'h0793; // 0x80001200
    mem[1153] <= 16'h14e3; // 0x80001204
    mem[1154] <= 16'h2717; // 0x80001208
    mem[1155] <= 16'h2703; // 0x8000120c
    mem[1156] <= 16'h0793; // 0x80001210
    mem[1157] <= 16'hda63; // 0x80001214
    mem[1158] <= 16'h2083; // 0x80001218
    mem[1159] <= 16'ha023; // 0x8000121c
    mem[1160] <= 16'h2403; // 0x80001220
    mem[1161] <= 16'h2483; // 0x80001224
    mem[1162] <= 16'h0113; // 0x80001228
    mem[1163] <= 16'h8067; // 0x8000122c
    mem[1164] <= 16'h2083; // 0x80001230
    mem[1165] <= 16'ha023; // 0x80001234
    mem[1166] <= 16'h2403; // 0x80001238
    mem[1167] <= 16'h2483; // 0x8000123c
    mem[1168] <= 16'h0113; // 0x80001240
    mem[1169] <= 16'h8067; // 0x80001244
    mem[1170] <= 16'h2083; // 0x80001248
    mem[1171] <= 16'h0793; // 0x8000124c
    mem[1172] <= 16'ha023; // 0x80001250
    mem[1173] <= 16'h2403; // 0x80001254
    mem[1174] <= 16'h2483; // 0x80001258
    mem[1175] <= 16'h0113; // 0x8000125c
    mem[1176] <= 16'h8067; // 0x80001260
    mem[1177] <= 16'h2717; // 0x80001264
    mem[1178] <= 16'h4703; // 0x80001268
    mem[1179] <= 16'h0793; // 0x8000126c
    mem[1180] <= 16'h0463; // 0x80001270
    mem[1181] <= 16'h8067; // 0x80001274
    mem[1182] <= 16'h2783; // 0x80001278
    mem[1183] <= 16'h2717; // 0x8000127c
    mem[1184] <= 16'h2703; // 0x80001280
    mem[1185] <= 16'h8793; // 0x80001284
    mem[1186] <= 16'h87b3; // 0x80001288
    mem[1187] <= 16'h2023; // 0x8000128c
    mem[1188] <= 16'h8067; // 0x80001290
    mem[1189] <= 16'h2617; // 0x80001294
    mem[1190] <= 16'h2603; // 0x80001298
    mem[1191] <= 16'h0a63; // 0x8000129c
    mem[1192] <= 16'h2783; // 0x800012a0
    mem[1193] <= 16'h2023; // 0x800012a4
    mem[1194] <= 16'h2617; // 0x800012a8
    mem[1195] <= 16'h2603; // 0x800012ac
    mem[1196] <= 16'h0613; // 0x800012b0
    mem[1197] <= 16'h2597; // 0x800012b4
    mem[1198] <= 16'ha583; // 0x800012b8
    mem[1199] <= 16'h0513; // 0x800012bc
    mem[1200] <= 16'hf06f; // 0x800012c0
    mem[1201] <= 16'h2797; // 0x800012c4
    mem[1202] <= 16'ha783; // 0x800012c8
    mem[1203] <= 16'h0113; // 0x800012cc
    mem[1204] <= 16'ha683; // 0x800012d0
    mem[1205] <= 16'h2423; // 0x800012d4
    mem[1206] <= 16'h2403; // 0x800012d8
    mem[1207] <= 16'h2623; // 0x800012dc
    mem[1208] <= 16'h2223; // 0x800012e0
    mem[1209] <= 16'h2023; // 0x800012e4
    mem[1210] <= 16'ha683; // 0x800012e8
    mem[1211] <= 16'h0493; // 0x800012ec
    mem[1212] <= 16'h0713; // 0x800012f0
    mem[1213] <= 16'h2223; // 0x800012f4
    mem[1214] <= 16'ha683; // 0x800012f8
    mem[1215] <= 16'h0513; // 0x800012fc
    mem[1216] <= 16'h2423; // 0x80001300
    mem[1217] <= 16'ha683; // 0x80001304
    mem[1218] <= 16'h2623; // 0x80001308
    mem[1219] <= 16'ha683; // 0x8000130c
    mem[1220] <= 16'h2823; // 0x80001310
    mem[1221] <= 16'ha683; // 0x80001314
    mem[1222] <= 16'h2a23; // 0x80001318
    mem[1223] <= 16'ha683; // 0x8000131c
    mem[1224] <= 16'h2c23; // 0x80001320
    mem[1225] <= 16'ha683; // 0x80001324
    mem[1226] <= 16'h2e23; // 0x80001328
    mem[1227] <= 16'ha683; // 0x8000132c
    mem[1228] <= 16'h2023; // 0x80001330
    mem[1229] <= 16'ha683; // 0x80001334
    mem[1230] <= 16'h2223; // 0x80001338
    mem[1231] <= 16'ha683; // 0x8000133c
    mem[1232] <= 16'h2423; // 0x80001340
    mem[1233] <= 16'ha783; // 0x80001344
    mem[1234] <= 16'h2623; // 0x80001348
    mem[1235] <= 16'ha623; // 0x8000134c
    mem[1236] <= 16'h2623; // 0x80001350
    mem[1237] <= 16'ha783; // 0x80001354
    mem[1238] <= 16'h2023; // 0x80001358
    mem[1239] <= 16'hf0ef; // 0x8000135c
    mem[1240] <= 16'h2783; // 0x80001360
    mem[1241] <= 16'h8e63; // 0x80001364
    mem[1242] <= 16'ha783; // 0x80001368
    mem[1243] <= 16'h2083; // 0x8000136c
    mem[1244] <= 16'h2403; // 0x80001370
    mem[1245] <= 16'ha703; // 0x80001374
    mem[1246] <= 16'ha023; // 0x80001378
    mem[1247] <= 16'ha703; // 0x8000137c
    mem[1248] <= 16'ha223; // 0x80001380
    mem[1249] <= 16'ha703; // 0x80001384
    mem[1250] <= 16'ha423; // 0x80001388
    mem[1251] <= 16'ha703; // 0x8000138c
    mem[1252] <= 16'ha623; // 0x80001390
    mem[1253] <= 16'ha703; // 0x80001394
    mem[1254] <= 16'ha823; // 0x80001398
    mem[1255] <= 16'ha703; // 0x8000139c
    mem[1256] <= 16'haa23; // 0x800013a0
    mem[1257] <= 16'ha703; // 0x800013a4
    mem[1258] <= 16'hac23; // 0x800013a8
    mem[1259] <= 16'ha703; // 0x800013ac
    mem[1260] <= 16'hae23; // 0x800013b0
    mem[1261] <= 16'ha703; // 0x800013b4
    mem[1262] <= 16'ha023; // 0x800013b8
    mem[1263] <= 16'ha703; // 0x800013bc
    mem[1264] <= 16'ha223; // 0x800013c0
    mem[1265] <= 16'ha703; // 0x800013c4
    mem[1266] <= 16'ha423; // 0x800013c8
    mem[1267] <= 16'ha783; // 0x800013cc
    mem[1268] <= 16'ha623; // 0x800013d0
    mem[1269] <= 16'h2483; // 0x800013d4
    mem[1270] <= 16'h0113; // 0x800013d8
    mem[1271] <= 16'h8067; // 0x800013dc
    mem[1272] <= 16'h0793; // 0x800013e0
    mem[1273] <= 16'h2623; // 0x800013e4
    mem[1274] <= 16'ha503; // 0x800013e8
    mem[1275] <= 16'h0593; // 0x800013ec
    mem[1276] <= 16'hf0ef; // 0x800013f0
    mem[1277] <= 16'h2797; // 0x800013f4
    mem[1278] <= 16'ha783; // 0x800013f8
    mem[1279] <= 16'ha783; // 0x800013fc
    mem[1280] <= 16'h2503; // 0x80001400
    mem[1281] <= 16'h0613; // 0x80001404
    mem[1282] <= 16'h2023; // 0x80001408
    mem[1283] <= 16'h2083; // 0x8000140c
    mem[1284] <= 16'h2403; // 0x80001410
    mem[1285] <= 16'h2483; // 0x80001414
    mem[1286] <= 16'h0593; // 0x80001418
    mem[1287] <= 16'h0113; // 0x8000141c
    mem[1288] <= 16'hf06f; // 0x80001420
    mem[1289] <= 16'h2717; // 0x80001424
    mem[1290] <= 16'h0713; // 0x80001428
    mem[1291] <= 16'h2683; // 0x8000142c
    mem[1292] <= 16'h2797; // 0x80001430
    mem[1293] <= 16'hc783; // 0x80001434
    mem[1294] <= 16'h8793; // 0x80001438
    mem[1295] <= 16'hb793; // 0x8000143c
    mem[1296] <= 16'he7b3; // 0x80001440
    mem[1297] <= 16'h2023; // 0x80001444
    mem[1298] <= 16'h0793; // 0x80001448
    mem[1299] <= 16'h2297; // 0x8000144c
    mem[1300] <= 16'h8c23; // 0x80001450
    mem[1301] <= 16'h8067; // 0x80001454
    mem[1302] <= 16'h0793; // 0x80001458
    mem[1303] <= 16'h2297; // 0x8000145c
    mem[1304] <= 16'h84a3; // 0x80001460
    mem[1305] <= 16'h2297; // 0x80001464
    mem[1306] <= 16'ha223; // 0x80001468
    mem[1307] <= 16'h8067; // 0x8000146c
    mem[1308] <= 16'h1737; // 0x80001470
    mem[1309] <= 16'h2783; // 0x80001474
    mem[1310] <= 16'hcee3; // 0x80001478
    mem[1311] <= 16'h7513; // 0x8000147c
    mem[1312] <= 16'h2023; // 0x80001480
    mem[1313] <= 16'h1737; // 0x80001484
    mem[1314] <= 16'h2783; // 0x80001488
    mem[1315] <= 16'hcee3; // 0x8000148c
    mem[1316] <= 16'h0513; // 0x80001490
    mem[1317] <= 16'h8067; // 0x80001494
    mem[1318] <= 16'h0793; // 0x80001498
    mem[1319] <= 16'h0713; // 0x8000149c
    mem[1320] <= 16'hca63; // 0x800014a0
    mem[1321] <= 16'h2783; // 0x800014a4
    mem[1322] <= 16'h9c63; // 0x800014a8
    mem[1323] <= 16'ha503; // 0x800014ac
    mem[1324] <= 16'h8793; // 0x800014b0
    mem[1325] <= 16'h0593; // 0x800014b4
    mem[1326] <= 16'h2023; // 0x800014b8
    mem[1327] <= 16'h8067; // 0x800014bc
    mem[1328] <= 16'h8693; // 0x800014c0
    mem[1329] <= 16'h2023; // 0x800014c4
    mem[1330] <= 16'h0593; // 0x800014c8
    mem[1331] <= 16'ha503; // 0x800014cc
    mem[1332] <= 16'h8067; // 0x800014d0
    mem[1333] <= 16'h2783; // 0x800014d4
    mem[1334] <= 16'h8793; // 0x800014d8
    mem[1335] <= 16'hf793; // 0x800014dc
    mem[1336] <= 16'h8693; // 0x800014e0
    mem[1337] <= 16'h2023; // 0x800014e4
    mem[1338] <= 16'ha583; // 0x800014e8
    mem[1339] <= 16'ha503; // 0x800014ec
    mem[1340] <= 16'h8067; // 0x800014f0
    mem[1341] <= 16'h0793; // 0x800014f4
    mem[1342] <= 16'h0713; // 0x800014f8
    mem[1343] <= 16'hce63; // 0x800014fc
    mem[1344] <= 16'h2783; // 0x80001500
    mem[1345] <= 16'ha503; // 0x80001504
    mem[1346] <= 16'h8793; // 0x80001508
    mem[1347] <= 16'h2023; // 0x8000150c
    mem[1348] <= 16'h5593; // 0x80001510
    mem[1349] <= 16'h8067; // 0x80001514
    mem[1350] <= 16'h2783; // 0x80001518
    mem[1351] <= 16'h8793; // 0x8000151c
    mem[1352] <= 16'hf793; // 0x80001520
    mem[1353] <= 16'h8693; // 0x80001524
    mem[1354] <= 16'h2023; // 0x80001528
    mem[1355] <= 16'ha583; // 0x8000152c
    mem[1356] <= 16'ha503; // 0x80001530
    mem[1357] <= 16'h8067; // 0x80001534
    mem[1358] <= 16'ha783; // 0x80001538
    mem[1359] <= 16'h8023; // 0x8000153c
    mem[1360] <= 16'ha783; // 0x80001540
    mem[1361] <= 16'h8793; // 0x80001544
    mem[1362] <= 16'ha023; // 0x80001548
    mem[1363] <= 16'h8067; // 0x8000154c
    mem[1364] <= 16'h0113; // 0x80001550
    mem[1365] <= 16'h2423; // 0x80001554
    mem[1366] <= 16'h8c13; // 0x80001558
    mem[1367] <= 16'h0693; // 0x8000155c
    mem[1368] <= 16'h2423; // 0x80001560
    mem[1369] <= 16'h2023; // 0x80001564
    mem[1370] <= 16'h2a23; // 0x80001568
    mem[1371] <= 16'h2823; // 0x8000156c
    mem[1372] <= 16'h2623; // 0x80001570
    mem[1373] <= 16'h2623; // 0x80001574
    mem[1374] <= 16'h2223; // 0x80001578
    mem[1375] <= 16'h2e23; // 0x8000157c
    mem[1376] <= 16'h2c23; // 0x80001580
    mem[1377] <= 16'h0913; // 0x80001584
    mem[1378] <= 16'h8413; // 0x80001588
    mem[1379] <= 16'h0a93; // 0x8000158c
    mem[1380] <= 16'h0b93; // 0x80001590
    mem[1381] <= 16'h10ef; // 0x80001594
    mem[1382] <= 16'h2023; // 0x80001598
    mem[1383] <= 16'h0b13; // 0x8000159c
    mem[1384] <= 16'h0263; // 0x800015a0
    mem[1385] <= 16'h0993; // 0x800015a4
    mem[1386] <= 16'h0493; // 0x800015a8
    mem[1387] <= 16'h8613; // 0x800015ac
    mem[1388] <= 16'h0693; // 0x800015b0
    mem[1389] <= 16'h0513; // 0x800015b4
    mem[1390] <= 16'h0593; // 0x800015b8
    mem[1391] <= 16'h10ef; // 0x800015bc
    mem[1392] <= 16'h8613; // 0x800015c0
    mem[1393] <= 16'h0693; // 0x800015c4
    mem[1394] <= 16'h0913; // 0x800015c8
    mem[1395] <= 16'h8413; // 0x800015cc
    mem[1396] <= 16'h10ef; // 0x800015d0
    mem[1397] <= 16'ha023; // 0x800015d4
    mem[1398] <= 16'h8a13; // 0x800015d8
    mem[1399] <= 16'h8993; // 0x800015dc
    mem[1400] <= 16'h0663; // 0x800015e0
    mem[1401] <= 16'h0493; // 0x800015e4
    mem[1402] <= 16'hf06f; // 0x800015e8
    mem[1403] <= 16'h7ce3; // 0x800015ec
    mem[1404] <= 16'h0413; // 0x800015f0
    mem[1405] <= 16'h5063; // 0x800015f4
    mem[1406] <= 16'h0593; // 0x800015f8
    mem[1407] <= 16'h8513; // 0x800015fc
    mem[1408] <= 16'h0413; // 0x80001600
    mem[1409] <= 16'hf0ef; // 0x80001604
    mem[1410] <= 16'h0793; // 0x80001608
    mem[1411] <= 16'h46e3; // 0x8000160c
    mem[1412] <= 16'h5263; // 0x80001610
    mem[1413] <= 16'h9413; // 0x80001614
    mem[1414] <= 16'h0433; // 0x80001618
    mem[1415] <= 16'h0993; // 0x8000161c
    mem[1416] <= 16'h0913; // 0x80001620
    mem[1417] <= 16'h0a13; // 0x80001624
    mem[1418] <= 16'h2783; // 0x80001628
    mem[1419] <= 16'h0593; // 0x8000162c
    mem[1420] <= 16'h8493; // 0x80001630
    mem[1421] <= 16'h0513; // 0x80001634
    mem[1422] <= 16'hf463; // 0x80001638
    mem[1423] <= 16'h0513; // 0x8000163c
    mem[1424] <= 16'h8533; // 0x80001640
    mem[1425] <= 16'hf0ef; // 0x80001644
    mem[1426] <= 16'h8793; // 0x80001648
    mem[1427] <= 16'h0413; // 0x8000164c
    mem[1428] <= 16'h4ce3; // 0x80001650
    mem[1429] <= 16'h2083; // 0x80001654
    mem[1430] <= 16'h2403; // 0x80001658
    mem[1431] <= 16'h2483; // 0x8000165c
    mem[1432] <= 16'h2903; // 0x80001660
    mem[1433] <= 16'h2983; // 0x80001664
    mem[1434] <= 16'h2a03; // 0x80001668
    mem[1435] <= 16'h2a83; // 0x8000166c
    mem[1436] <= 16'h2b03; // 0x80001670
    mem[1437] <= 16'h2b83; // 0x80001674
    mem[1438] <= 16'h2c03; // 0x80001678
    mem[1439] <= 16'h0113; // 0x8000167c
    mem[1440] <= 16'h8067; // 0x80001680
    mem[1441] <= 16'h70e3; // 0x80001684
    mem[1442] <= 16'h0a13; // 0x80001688
    mem[1443] <= 16'h0413; // 0x8000168c
    mem[1444] <= 16'h0493; // 0x80001690
    mem[1445] <= 16'h42e3; // 0x80001694
    mem[1446] <= 16'hf06f; // 0x80001698
    mem[1447] <= 16'h0113; // 0x8000169c
    mem[1448] <= 16'h2423; // 0x800016a0
    mem[1449] <= 16'h2023; // 0x800016a4
    mem[1450] <= 16'h8413; // 0x800016a8
    mem[1451] <= 16'h0913; // 0x800016ac
    mem[1452] <= 16'h2c23; // 0x800016b0
    mem[1453] <= 16'h0613; // 0x800016b4
    mem[1454] <= 16'h0a13; // 0x800016b8
    mem[1455] <= 16'h0693; // 0x800016bc
    mem[1456] <= 16'h0513; // 0x800016c0
    mem[1457] <= 16'h0593; // 0x800016c4
    mem[1458] <= 16'h2823; // 0x800016c8
    mem[1459] <= 16'h2623; // 0x800016cc
    mem[1460] <= 16'h2423; // 0x800016d0
    mem[1461] <= 16'h2223; // 0x800016d4
    mem[1462] <= 16'h2623; // 0x800016d8
    mem[1463] <= 16'h2223; // 0x800016dc
    mem[1464] <= 16'h2e23; // 0x800016e0
    mem[1465] <= 16'h2a23; // 0x800016e4
    mem[1466] <= 16'h0b13; // 0x800016e8
    mem[1467] <= 16'h8c93; // 0x800016ec
    mem[1468] <= 16'h0c13; // 0x800016f0
    mem[1469] <= 16'h10ef; // 0x800016f4
    mem[1470] <= 16'h2023; // 0x800016f8
    mem[1471] <= 16'h0b93; // 0x800016fc
    mem[1472] <= 16'h0463; // 0x80001700
    mem[1473] <= 16'h0993; // 0x80001704
    mem[1474] <= 16'h0493; // 0x80001708
    mem[1475] <= 16'h0613; // 0x8000170c
    mem[1476] <= 16'h0693; // 0x80001710
    mem[1477] <= 16'h0513; // 0x80001714
    mem[1478] <= 16'h0593; // 0x80001718
    mem[1479] <= 16'h10ef; // 0x8000171c
    mem[1480] <= 16'h0613; // 0x80001720
    mem[1481] <= 16'h0693; // 0x80001724
    mem[1482] <= 16'h0913; // 0x80001728
    mem[1483] <= 16'h8413; // 0x8000172c
    mem[1484] <= 16'h10ef; // 0x80001730
    mem[1485] <= 16'ha023; // 0x80001734
    mem[1486] <= 16'h8a93; // 0x80001738
    mem[1487] <= 16'h8993; // 0x8000173c
    mem[1488] <= 16'h8663; // 0x80001740
    mem[1489] <= 16'h8493; // 0x80001744
    mem[1490] <= 16'hf06f; // 0x80001748
    mem[1491] <= 16'h7ce3; // 0x8000174c
    mem[1492] <= 16'h8413; // 0x80001750
    mem[1493] <= 16'hd063; // 0x80001754
    mem[1494] <= 16'h0593; // 0x80001758
    mem[1495] <= 16'h0513; // 0x8000175c
    mem[1496] <= 16'h0413; // 0x80001760
    mem[1497] <= 16'hf0ef; // 0x80001764
    mem[1498] <= 16'h0793; // 0x80001768
    mem[1499] <= 16'hc6e3; // 0x8000176c
    mem[1500] <= 16'h5263; // 0x80001770
    mem[1501] <= 16'h9413; // 0x80001774
    mem[1502] <= 16'h0433; // 0x80001778
    mem[1503] <= 16'h0993; // 0x8000177c
    mem[1504] <= 16'h0913; // 0x80001780
    mem[1505] <= 16'h0a93; // 0x80001784
    mem[1506] <= 16'h2783; // 0x80001788
    mem[1507] <= 16'h0593; // 0x8000178c
    mem[1508] <= 16'h8493; // 0x80001790
    mem[1509] <= 16'h0513; // 0x80001794
    mem[1510] <= 16'hf463; // 0x80001798
    mem[1511] <= 16'h8513; // 0x8000179c
    mem[1512] <= 16'h8533; // 0x800017a0
    mem[1513] <= 16'hf0ef; // 0x800017a4
    mem[1514] <= 16'h8793; // 0x800017a8
    mem[1515] <= 16'h0413; // 0x800017ac
    mem[1516] <= 16'h4ce3; // 0x800017b0
    mem[1517] <= 16'h2083; // 0x800017b4
    mem[1518] <= 16'h2403; // 0x800017b8
    mem[1519] <= 16'h2483; // 0x800017bc
    mem[1520] <= 16'h2903; // 0x800017c0
    mem[1521] <= 16'h2983; // 0x800017c4
    mem[1522] <= 16'h2a03; // 0x800017c8
    mem[1523] <= 16'h2a83; // 0x800017cc
    mem[1524] <= 16'h2b03; // 0x800017d0
    mem[1525] <= 16'h2b83; // 0x800017d4
    mem[1526] <= 16'h2c03; // 0x800017d8
    mem[1527] <= 16'h2c83; // 0x800017dc
    mem[1528] <= 16'h0113; // 0x800017e0
    mem[1529] <= 16'h8067; // 0x800017e4
    mem[1530] <= 16'h7ee3; // 0x800017e8
    mem[1531] <= 16'h0a93; // 0x800017ec
    mem[1532] <= 16'h8413; // 0x800017f0
    mem[1533] <= 16'h0493; // 0x800017f4
    mem[1534] <= 16'hc0e3; // 0x800017f8
    mem[1535] <= 16'hf06f; // 0x800017fc
    mem[1536] <= 16'h27f3; // 0x80001800
    mem[1537] <= 16'h1063; // 0x80001804
    mem[1538] <= 16'h2717; // 0x80001808
    mem[1539] <= 16'h2703; // 0x8000180c
    mem[1540] <= 16'h87b3; // 0x80001810
    mem[1541] <= 16'h2717; // 0x80001814
    mem[1542] <= 16'h0713; // 0x80001818
    mem[1543] <= 16'h2297; // 0x8000181c
    mem[1544] <= 16'hae23; // 0x80001820
    mem[1545] <= 16'h2717; // 0x80001824
    mem[1546] <= 16'h0713; // 0x80001828
    mem[1547] <= 16'h2023; // 0x8000182c
    mem[1548] <= 16'h27f3; // 0x80001830
    mem[1549] <= 16'h1063; // 0x80001834
    mem[1550] <= 16'h2697; // 0x80001838
    mem[1551] <= 16'ha683; // 0x8000183c
    mem[1552] <= 16'h87b3; // 0x80001840
    mem[1553] <= 16'h2697; // 0x80001844
    mem[1554] <= 16'h8693; // 0x80001848
    mem[1555] <= 16'h2297; // 0x8000184c
    mem[1556] <= 16'ha823; // 0x80001850
    mem[1557] <= 16'h2223; // 0x80001854
    mem[1558] <= 16'h8067; // 0x80001858
    mem[1559] <= 16'h1513; // 0x8000185c
    mem[1560] <= 16'hf697; // 0x80001860
    mem[1561] <= 16'h8693; // 0x80001864
    mem[1562] <= 16'h6713; // 0x80001868
    mem[1563] <= 16'h0793; // 0x8000186c
    mem[1564] <= 16'ha023; // 0x80001870
    mem[1565] <= 16'ha223; // 0x80001874
    mem[1566] <= 16'h006f; // 0x80001878
    mem[1567] <= 16'h0113; // 0x8000187c
    mem[1568] <= 16'h0513; // 0x80001880
    mem[1569] <= 16'h2623; // 0x80001884
    mem[1570] <= 16'hf0ef; // 0x80001888
    mem[1571] <= 16'h0113; // 0x8000188c
    mem[1572] <= 16'h2623; // 0x80001890
    mem[1573] <= 16'hf0ef; // 0x80001894
    mem[1574] <= 16'h0113; // 0x80001898
    mem[1575] <= 16'h0513; // 0x8000189c
    mem[1576] <= 16'h2623; // 0x800018a0
    mem[1577] <= 16'hf0ef; // 0x800018a4
    mem[1578] <= 16'h0463; // 0x800018a8
    mem[1579] <= 16'h006f; // 0x800018ac
    mem[1580] <= 16'h8067; // 0x800018b0
    mem[1581] <= 16'he7b3; // 0x800018b4
    mem[1582] <= 16'he7b3; // 0x800018b8
    mem[1583] <= 16'hf793; // 0x800018bc
    mem[1584] <= 16'h8863; // 0x800018c0
    mem[1585] <= 16'h0833; // 0x800018c4
    mem[1586] <= 16'h7663; // 0x800018c8
    mem[1587] <= 16'h8713; // 0x800018cc
    mem[1588] <= 16'h0693; // 0x800018d0
    mem[1589] <= 16'h3733; // 0x800018d4
    mem[1590] <= 16'hb6b3; // 0x800018d8
    mem[1591] <= 16'h67b3; // 0x800018dc
    mem[1592] <= 16'h4713; // 0x800018e0
    mem[1593] <= 16'hc693; // 0x800018e4
    mem[1594] <= 16'hf793; // 0x800018e8
    mem[1595] <= 16'h6733; // 0x800018ec
    mem[1596] <= 16'hb793; // 0x800018f0
    mem[1597] <= 16'hf7b3; // 0x800018f4
    mem[1598] <= 16'h8e63; // 0x800018f8
    mem[1599] <= 16'h3793; // 0x800018fc
    mem[1600] <= 16'h9a63; // 0x80001900
    mem[1601] <= 16'h0793; // 0x80001904
    mem[1602] <= 16'hd793; // 0x80001908
    mem[1603] <= 16'h8793; // 0x8000190c
    mem[1604] <= 16'h9313; // 0x80001910
    mem[1605] <= 16'h0893; // 0x80001914
    mem[1606] <= 16'h8693; // 0x80001918
    mem[1607] <= 16'h0713; // 0x8000191c
    mem[1608] <= 16'hae03; // 0x80001920
    mem[1609] <= 16'h0713; // 0x80001924
    mem[1610] <= 16'h8693; // 0x80001928
    mem[1611] <= 16'ha023; // 0x8000192c
    mem[1612] <= 16'h8893; // 0x80001930
    mem[1613] <= 16'h66e3; // 0x80001934
    mem[1614] <= 16'h85b3; // 0x80001938
    mem[1615] <= 16'h07b3; // 0x8000193c
    mem[1616] <= 16'h0663; // 0x80001940
    mem[1617] <= 16'hc683; // 0x80001944
    mem[1618] <= 16'h8713; // 0x80001948
    mem[1619] <= 16'h8023; // 0x8000194c
    mem[1620] <= 16'h7e63; // 0x80001950
    mem[1621] <= 16'hc683; // 0x80001954
    mem[1622] <= 16'h8713; // 0x80001958
    mem[1623] <= 16'h80a3; // 0x8000195c
    mem[1624] <= 16'h7863; // 0x80001960
    mem[1625] <= 16'hc703; // 0x80001964
    mem[1626] <= 16'h8123; // 0x80001968
    mem[1627] <= 16'h8067; // 0x8000196c
    mem[1628] <= 16'h0633; // 0x80001970
    mem[1629] <= 16'h7c63; // 0x80001974
    mem[1630] <= 16'h0793; // 0x80001978
    mem[1631] <= 16'h8593; // 0x8000197c
    mem[1632] <= 16'ha703; // 0x80001980
    mem[1633] <= 16'h8793; // 0x80001984
    mem[1634] <= 16'hae23; // 0x80001988
    mem[1635] <= 16'he8e3; // 0x8000198c
    mem[1636] <= 16'h8067; // 0x80001990
    mem[1637] <= 16'h0793; // 0x80001994
    mem[1638] <= 16'h8593; // 0x80001998
    mem[1639] <= 16'hc703; // 0x8000199c
    mem[1640] <= 16'h8793; // 0x800019a0
    mem[1641] <= 16'h8fa3; // 0x800019a4
    mem[1642] <= 16'h18e3; // 0x800019a8
    mem[1643] <= 16'h8067; // 0x800019ac
    mem[1644] <= 16'h8067; // 0x800019b0
    mem[1645] <= 16'h8067; // 0x800019b4
    mem[1646] <= 16'h0113; // 0x800019b8
    mem[1647] <= 16'h67b3; // 0x800019bc
    mem[1648] <= 16'h2423; // 0x800019c0
    mem[1649] <= 16'h2623; // 0x800019c4
    mem[1650] <= 16'hf793; // 0x800019c8
    mem[1651] <= 16'h0413; // 0x800019cc
    mem[1652] <= 16'h8663; // 0x800019d0
    mem[1653] <= 16'h0633; // 0x800019d4
    mem[1654] <= 16'h7863; // 0x800019d8
    mem[1655] <= 16'h0633; // 0x800019dc
    mem[1656] <= 16'hf593; // 0x800019e0
    mem[1657] <= 16'hf0ef; // 0x800019e4
    mem[1658] <= 16'h2083; // 0x800019e8
    mem[1659] <= 16'h0513; // 0x800019ec
    mem[1660] <= 16'h2403; // 0x800019f0
    mem[1661] <= 16'h0113; // 0x800019f4
    mem[1662] <= 16'h8067; // 0x800019f8
    mem[1663] <= 16'hf713; // 0x800019fc
    mem[1664] <= 16'h1593; // 0x80001a00
    mem[1665] <= 16'h6733; // 0x80001a04
    mem[1666] <= 16'h1793; // 0x80001a08
    mem[1667] <= 16'h0633; // 0x80001a0c
    mem[1668] <= 16'h6733; // 0x80001a10
    mem[1669] <= 16'h7ae3; // 0x80001a14
    mem[1670] <= 16'h0793; // 0x80001a18
    mem[1671] <= 16'h8793; // 0x80001a1c
    mem[1672] <= 16'hae23; // 0x80001a20
    mem[1673] <= 16'hece3; // 0x80001a24
    mem[1674] <= 16'h2083; // 0x80001a28
    mem[1675] <= 16'h0513; // 0x80001a2c
    mem[1676] <= 16'h2403; // 0x80001a30
    mem[1677] <= 16'h0113; // 0x80001a34
    mem[1678] <= 16'h8067; // 0x80001a38
    mem[1679] <= 16'h0113; // 0x80001a3c
    mem[1680] <= 16'h2423; // 0x80001a40
    mem[1681] <= 16'h2223; // 0x80001a44
    mem[1682] <= 16'h0493; // 0x80001a48
    mem[1683] <= 16'h0413; // 0x80001a4c
    mem[1684] <= 16'h8433; // 0x80001a50
    mem[1685] <= 16'h0613; // 0x80001a54
    mem[1686] <= 16'h4597; // 0x80001a58
    mem[1687] <= 16'h8593; // 0x80001a5c
    mem[1688] <= 16'h0513; // 0x80001a60
    mem[1689] <= 16'h2623; // 0x80001a64
    mem[1690] <= 16'h2023; // 0x80001a68
    mem[1691] <= 16'h0913; // 0x80001a6c
    mem[1692] <= 16'hf0ef; // 0x80001a70
    mem[1693] <= 16'h0613; // 0x80001a74
    mem[1694] <= 16'h0533; // 0x80001a78
    mem[1695] <= 16'h0633; // 0x80001a7c
    mem[1696] <= 16'h2083; // 0x80001a80
    mem[1697] <= 16'h2403; // 0x80001a84
    mem[1698] <= 16'h2483; // 0x80001a88
    mem[1699] <= 16'h2903; // 0x80001a8c
    mem[1700] <= 16'h0593; // 0x80001a90
    mem[1701] <= 16'h0113; // 0x80001a94
    mem[1702] <= 16'hf06f; // 0x80001a98
    mem[1703] <= 16'h4783; // 0x80001a9c
    mem[1704] <= 16'h8e63; // 0x80001aa0
    mem[1705] <= 16'h0793; // 0x80001aa4
    mem[1706] <= 16'h8793; // 0x80001aa8
    mem[1707] <= 16'hc703; // 0x80001aac
    mem[1708] <= 16'h1ce3; // 0x80001ab0
    mem[1709] <= 16'h8533; // 0x80001ab4
    mem[1710] <= 16'h8067; // 0x80001ab8
    mem[1711] <= 16'h0513; // 0x80001abc
    mem[1712] <= 16'h8067; // 0x80001ac0
    mem[1713] <= 16'h0113; // 0x80001ac4
    mem[1714] <= 16'h2623; // 0x80001ac8
    mem[1715] <= 16'h0993; // 0x80001acc
    mem[1716] <= 16'h2823; // 0x80001ad0
    mem[1717] <= 16'h0913; // 0x80001ad4
    mem[1718] <= 16'h8513; // 0x80001ad8
    mem[1719] <= 16'h2c23; // 0x80001adc
    mem[1720] <= 16'h2a23; // 0x80001ae0
    mem[1721] <= 16'h2e23; // 0x80001ae4
    mem[1722] <= 16'h0493; // 0x80001ae8
    mem[1723] <= 16'h1437; // 0x80001aec
    mem[1724] <= 16'hf0ef; // 0x80001af0
    mem[1725] <= 16'hf863; // 0x80001af4
    mem[1726] <= 16'h2783; // 0x80001af8
    mem[1727] <= 16'hcee3; // 0x80001afc
    mem[1728] <= 16'h4783; // 0x80001b00
    mem[1729] <= 16'h2023; // 0x80001b04
    mem[1730] <= 16'h2783; // 0x80001b08
    mem[1731] <= 16'hcee3; // 0x80001b0c
    mem[1732] <= 16'h8513; // 0x80001b10
    mem[1733] <= 16'h8493; // 0x80001b14
    mem[1734] <= 16'h0913; // 0x80001b18
    mem[1735] <= 16'hf0ef; // 0x80001b1c
    mem[1736] <= 16'hece3; // 0x80001b20
    mem[1737] <= 16'h2083; // 0x80001b24
    mem[1738] <= 16'h2403; // 0x80001b28
    mem[1739] <= 16'h2483; // 0x80001b2c
    mem[1740] <= 16'h2903; // 0x80001b30
    mem[1741] <= 16'h2983; // 0x80001b34
    mem[1742] <= 16'h0113; // 0x80001b38
    mem[1743] <= 16'h8067; // 0x80001b3c
    mem[1744] <= 16'h0113; // 0x80001b40
    mem[1745] <= 16'h2623; // 0x80001b44
    mem[1746] <= 16'h7793; // 0x80001b48
    mem[1747] <= 16'h0693; // 0x80001b4c
    mem[1748] <= 16'h0713; // 0x80001b50
    mem[1749] <= 16'hf463; // 0x80001b54
    mem[1750] <= 16'h0713; // 0x80001b58
    mem[1751] <= 16'h8733; // 0x80001b5c
    mem[1752] <= 16'h5793; // 0x80001b60
    mem[1753] <= 16'h0da3; // 0x80001b64
    mem[1754] <= 16'hf793; // 0x80001b68
    mem[1755] <= 16'h0693; // 0x80001b6c
    mem[1756] <= 16'h0713; // 0x80001b70
    mem[1757] <= 16'he463; // 0x80001b74
    mem[1758] <= 16'h0713; // 0x80001b78
    mem[1759] <= 16'h8733; // 0x80001b7c
    mem[1760] <= 16'h5793; // 0x80001b80
    mem[1761] <= 16'h0d23; // 0x80001b84
    mem[1762] <= 16'hf793; // 0x80001b88
    mem[1763] <= 16'h0693; // 0x80001b8c
    mem[1764] <= 16'h0713; // 0x80001b90
    mem[1765] <= 16'he463; // 0x80001b94
    mem[1766] <= 16'h0713; // 0x80001b98
    mem[1767] <= 16'h8733; // 0x80001b9c
    mem[1768] <= 16'h5793; // 0x80001ba0
    mem[1769] <= 16'h0ca3; // 0x80001ba4
    mem[1770] <= 16'hf793; // 0x80001ba8
    mem[1771] <= 16'h0693; // 0x80001bac
    mem[1772] <= 16'h0713; // 0x80001bb0
    mem[1773] <= 16'he463; // 0x80001bb4
    mem[1774] <= 16'h0713; // 0x80001bb8
    mem[1775] <= 16'h8733; // 0x80001bbc
    mem[1776] <= 16'h5793; // 0x80001bc0
    mem[1777] <= 16'h0c23; // 0x80001bc4
    mem[1778] <= 16'hf793; // 0x80001bc8
    mem[1779] <= 16'h0693; // 0x80001bcc
    mem[1780] <= 16'h0713; // 0x80001bd0
    mem[1781] <= 16'he463; // 0x80001bd4
    mem[1782] <= 16'h0713; // 0x80001bd8
    mem[1783] <= 16'h8733; // 0x80001bdc
    mem[1784] <= 16'h5793; // 0x80001be0
    mem[1785] <= 16'h0ba3; // 0x80001be4
    mem[1786] <= 16'hf793; // 0x80001be8
    mem[1787] <= 16'h0693; // 0x80001bec
    mem[1788] <= 16'h0713; // 0x80001bf0
    mem[1789] <= 16'he463; // 0x80001bf4
    mem[1790] <= 16'h0713; // 0x80001bf8
    mem[1791] <= 16'h8733; // 0x80001bfc
    mem[1792] <= 16'h5793; // 0x80001c00
    mem[1793] <= 16'h0b23; // 0x80001c04
    mem[1794] <= 16'hf793; // 0x80001c08
    mem[1795] <= 16'h0693; // 0x80001c0c
    mem[1796] <= 16'h0713; // 0x80001c10
    mem[1797] <= 16'he463; // 0x80001c14
    mem[1798] <= 16'h0713; // 0x80001c18
    mem[1799] <= 16'h87b3; // 0x80001c1c
    mem[1800] <= 16'h0aa3; // 0x80001c20
    mem[1801] <= 16'h5513; // 0x80001c24
    mem[1802] <= 16'h0713; // 0x80001c28
    mem[1803] <= 16'h0793; // 0x80001c2c
    mem[1804] <= 16'h6463; // 0x80001c30
    mem[1805] <= 16'h0793; // 0x80001c34
    mem[1806] <= 16'h0533; // 0x80001c38
    mem[1807] <= 16'h0a23; // 0x80001c3c
    mem[1808] <= 16'hf793; // 0x80001c40
    mem[1809] <= 16'h0693; // 0x80001c44
    mem[1810] <= 16'h0713; // 0x80001c48
    mem[1811] <= 16'he463; // 0x80001c4c
    mem[1812] <= 16'h0713; // 0x80001c50
    mem[1813] <= 16'h8733; // 0x80001c54
    mem[1814] <= 16'hd793; // 0x80001c58
    mem[1815] <= 16'h09a3; // 0x80001c5c
    mem[1816] <= 16'hf793; // 0x80001c60
    mem[1817] <= 16'h0693; // 0x80001c64
    mem[1818] <= 16'h0713; // 0x80001c68
    mem[1819] <= 16'he463; // 0x80001c6c
    mem[1820] <= 16'h0713; // 0x80001c70
    mem[1821] <= 16'h8733; // 0x80001c74
    mem[1822] <= 16'hd793; // 0x80001c78
    mem[1823] <= 16'h0923; // 0x80001c7c
    mem[1824] <= 16'hf793; // 0x80001c80
    mem[1825] <= 16'h0693; // 0x80001c84
    mem[1826] <= 16'h0713; // 0x80001c88
    mem[1827] <= 16'he463; // 0x80001c8c
    mem[1828] <= 16'h0713; // 0x80001c90
    mem[1829] <= 16'h8733; // 0x80001c94
    mem[1830] <= 16'hd793; // 0x80001c98
    mem[1831] <= 16'h08a3; // 0x80001c9c
    mem[1832] <= 16'hf793; // 0x80001ca0
    mem[1833] <= 16'h0693; // 0x80001ca4
    mem[1834] <= 16'h0713; // 0x80001ca8
    mem[1835] <= 16'he463; // 0x80001cac
    mem[1836] <= 16'h0713; // 0x80001cb0
    mem[1837] <= 16'h8733; // 0x80001cb4
    mem[1838] <= 16'hd793; // 0x80001cb8
    mem[1839] <= 16'h0823; // 0x80001cbc
    mem[1840] <= 16'hf793; // 0x80001cc0
    mem[1841] <= 16'h0693; // 0x80001cc4
    mem[1842] <= 16'h0713; // 0x80001cc8
    mem[1843] <= 16'he463; // 0x80001ccc
    mem[1844] <= 16'h0713; // 0x80001cd0
    mem[1845] <= 16'h8733; // 0x80001cd4
    mem[1846] <= 16'hd793; // 0x80001cd8
    mem[1847] <= 16'h07a3; // 0x80001cdc
    mem[1848] <= 16'hf793; // 0x80001ce0
    mem[1849] <= 16'h0693; // 0x80001ce4
    mem[1850] <= 16'h0713; // 0x80001ce8
    mem[1851] <= 16'he463; // 0x80001cec
    mem[1852] <= 16'h0713; // 0x80001cf0
    mem[1853] <= 16'h8733; // 0x80001cf4
    mem[1854] <= 16'hd793; // 0x80001cf8
    mem[1855] <= 16'h0723; // 0x80001cfc
    mem[1856] <= 16'hf793; // 0x80001d00
    mem[1857] <= 16'h0693; // 0x80001d04
    mem[1858] <= 16'h0713; // 0x80001d08
    mem[1859] <= 16'he463; // 0x80001d0c
    mem[1860] <= 16'h0713; // 0x80001d10
    mem[1861] <= 16'h87b3; // 0x80001d14
    mem[1862] <= 16'h06a3; // 0x80001d18
    mem[1863] <= 16'hd593; // 0x80001d1c
    mem[1864] <= 16'h0713; // 0x80001d20
    mem[1865] <= 16'h0793; // 0x80001d24
    mem[1866] <= 16'h6463; // 0x80001d28
    mem[1867] <= 16'h0793; // 0x80001d2c
    mem[1868] <= 16'h85b3; // 0x80001d30
    mem[1869] <= 16'h0513; // 0x80001d34
    mem[1870] <= 16'h0623; // 0x80001d38
    mem[1871] <= 16'h0e23; // 0x80001d3c
    mem[1872] <= 16'hf0ef; // 0x80001d40
    mem[1873] <= 16'h2083; // 0x80001d44
    mem[1874] <= 16'h0113; // 0x80001d48
    mem[1875] <= 16'h8067; // 0x80001d4c
    mem[1876] <= 16'h8863; // 0x80001d50
    mem[1877] <= 16'h4783; // 0x80001d54
    mem[1878] <= 16'h8463; // 0x80001d58
    mem[1879] <= 16'h05b3; // 0x80001d5c
    mem[1880] <= 16'h0793; // 0x80001d60
    mem[1881] <= 16'h006f; // 0x80001d64
    mem[1882] <= 16'hc703; // 0x80001d68
    mem[1883] <= 16'h0663; // 0x80001d6c
    mem[1884] <= 16'h8793; // 0x80001d70
    mem[1885] <= 16'h9ae3; // 0x80001d74
    mem[1886] <= 16'h8533; // 0x80001d78
    mem[1887] <= 16'h8067; // 0x80001d7c
    mem[1888] <= 16'h0513; // 0x80001d80
    mem[1889] <= 16'h8067; // 0x80001d84
    mem[1890] <= 16'h0113; // 0x80001d88
    mem[1891] <= 16'h2c23; // 0x80001d8c
    mem[1892] <= 16'h2823; // 0x80001d90
    mem[1893] <= 16'h2623; // 0x80001d94
    mem[1894] <= 16'h2423; // 0x80001d98
    mem[1895] <= 16'h2223; // 0x80001d9c
    mem[1896] <= 16'h2023; // 0x80001da0
    mem[1897] <= 16'h2e23; // 0x80001da4
    mem[1898] <= 16'h2a23; // 0x80001da8
    mem[1899] <= 16'h2e23; // 0x80001dac
    mem[1900] <= 16'h2c23; // 0x80001db0
    mem[1901] <= 16'h2a23; // 0x80001db4
    mem[1902] <= 16'h2823; // 0x80001db8
    mem[1903] <= 16'h0913; // 0x80001dbc
    mem[1904] <= 16'h8413; // 0x80001dc0
    mem[1905] <= 16'h2623; // 0x80001dc4
    mem[1906] <= 16'h1997; // 0x80001dc8
    mem[1907] <= 16'h8993; // 0x80001dcc
    mem[1908] <= 16'h0b13; // 0x80001dd0
    mem[1909] <= 16'h0a93; // 0x80001dd4
    mem[1910] <= 16'h0a13; // 0x80001dd8
    mem[1911] <= 16'h4503; // 0x80001ddc
    mem[1912] <= 16'h0493; // 0x80001de0
    mem[1913] <= 16'h0e63; // 0x80001de4
    mem[1914] <= 16'h0863; // 0x80001de8
    mem[1915] <= 16'h0593; // 0x80001dec
    mem[1916] <= 16'h0413; // 0x80001df0
    mem[1917] <= 16'hf0ef; // 0x80001df4
    mem[1918] <= 16'h4503; // 0x80001df8
    mem[1919] <= 16'h16e3; // 0x80001dfc
    mem[1920] <= 16'h2603; // 0x80001e00
    mem[1921] <= 16'h4e03; // 0x80001e04
    mem[1922] <= 16'h0c93; // 0x80001e08
    mem[1923] <= 16'h0493; // 0x80001e0c
    mem[1924] <= 16'h0893; // 0x80001e10
    mem[1925] <= 16'h8793; // 0x80001e14
    mem[1926] <= 16'h0813; // 0x80001e18
    mem[1927] <= 16'h0b93; // 0x80001e1c
    mem[1928] <= 16'h8c13; // 0x80001e20
    mem[1929] <= 16'h0593; // 0x80001e24
    mem[1930] <= 16'h0693; // 0x80001e28
    mem[1931] <= 16'h0513; // 0x80001e2c
    mem[1932] <= 16'h0313; // 0x80001e30
    mem[1933] <= 16'h0713; // 0x80001e34
    mem[1934] <= 16'h7713; // 0x80001e38
    mem[1935] <= 16'h8413; // 0x80001e3c
    mem[1936] <= 16'he463; // 0x80001e40
    mem[1937] <= 16'h1713; // 0x80001e44
    mem[1938] <= 16'h0733; // 0x80001e48
    mem[1939] <= 16'h2703; // 0x80001e4c
    mem[1940] <= 16'h0733; // 0x80001e50
    mem[1941] <= 16'h0067; // 0x80001e54
    mem[1942] <= 16'h2083; // 0x80001e58
    mem[1943] <= 16'h2403; // 0x80001e5c
    mem[1944] <= 16'h2483; // 0x80001e60
    mem[1945] <= 16'h2903; // 0x80001e64
    mem[1946] <= 16'h2983; // 0x80001e68
    mem[1947] <= 16'h2a03; // 0x80001e6c
    mem[1948] <= 16'h2a83; // 0x80001e70
    mem[1949] <= 16'h2b03; // 0x80001e74
    mem[1950] <= 16'h2b83; // 0x80001e78
    mem[1951] <= 16'h2c03; // 0x80001e7c
    mem[1952] <= 16'h2c83; // 0x80001e80
    mem[1953] <= 16'h2d03; // 0x80001e84
    mem[1954] <= 16'h0113; // 0x80001e88
    mem[1955] <= 16'h8067; // 0x80001e8c
    mem[1956] <= 16'h5463; // 0x80001e90
    mem[1957] <= 16'h0c13; // 0x80001e94
    mem[1958] <= 16'hce03; // 0x80001e98
    mem[1959] <= 16'h0793; // 0x80001e9c
    mem[1960] <= 16'hf06f; // 0x80001ea0
    mem[1961] <= 16'h1c63; // 0x80001ea4
    mem[1962] <= 16'h0493; // 0x80001ea8
    mem[1963] <= 16'h0513; // 0x80001eac
    mem[1964] <= 16'hf0ef; // 0x80001eb0
    mem[1965] <= 16'h0613; // 0x80001eb4
    mem[1966] <= 16'h8693; // 0x80001eb8
    mem[1967] <= 16'h8813; // 0x80001ebc
    mem[1968] <= 16'h0793; // 0x80001ec0
    mem[1969] <= 16'h8713; // 0x80001ec4
    mem[1970] <= 16'h0513; // 0x80001ec8
    mem[1971] <= 16'hf0ef; // 0x80001ecc
    mem[1972] <= 16'hf06f; // 0x80001ed0
    mem[1973] <= 16'h1063; // 0x80001ed4
    mem[1974] <= 16'h0593; // 0x80001ed8
    mem[1975] <= 16'h0513; // 0x80001edc
    mem[1976] <= 16'hf0ef; // 0x80001ee0
    mem[1977] <= 16'hf06f; // 0x80001ee4
    mem[1978] <= 16'ha483; // 0x80001ee8
    mem[1979] <= 16'hce03; // 0x80001eec
    mem[1980] <= 16'h8893; // 0x80001ef0
    mem[1981] <= 16'h0793; // 0x80001ef4
    mem[1982] <= 16'h0813; // 0x80001ef8
    mem[1983] <= 16'h5ce3; // 0x80001efc
    mem[1984] <= 16'h8c13; // 0x80001f00
    mem[1985] <= 16'h0493; // 0x80001f04
    mem[1986] <= 16'hf06f; // 0x80001f08
    mem[1987] <= 16'hce03; // 0x80001f0c
    mem[1988] <= 16'h0b93; // 0x80001f10
    mem[1989] <= 16'h0793; // 0x80001f14
    mem[1990] <= 16'hf06f; // 0x80001f18
    mem[1991] <= 16'hce03; // 0x80001f1c
    mem[1992] <= 16'h8b93; // 0x80001f20
    mem[1993] <= 16'h0793; // 0x80001f24
    mem[1994] <= 16'hf06f; // 0x80001f28
    mem[1995] <= 16'hce83; // 0x80001f2c
    mem[1996] <= 16'h0493; // 0x80001f30
    mem[1997] <= 16'h8793; // 0x80001f34
    mem[1998] <= 16'h6863; // 0x80001f38
    mem[1999] <= 16'h0793; // 0x80001f3c
    mem[2000] <= 16'h9713; // 0x80001f40
    mem[2001] <= 16'h04b3; // 0x80001f44
    mem[2002] <= 16'h8793; // 0x80001f48
    mem[2003] <= 16'h9493; // 0x80001f4c
    mem[2004] <= 16'h84b3; // 0x80001f50
    mem[2005] <= 16'hce83; // 0x80001f54
    mem[2006] <= 16'h8493; // 0x80001f58
    mem[2007] <= 16'h8713; // 0x80001f5c
    mem[2008] <= 16'h70e3; // 0x80001f60
    mem[2009] <= 16'h8e13; // 0x80001f64
    mem[2010] <= 16'hf06f; // 0x80001f68
    mem[2011] <= 16'h1c63; // 0x80001f6c
    mem[2012] <= 16'h2503; // 0x80001f70
    mem[2013] <= 16'h0593; // 0x80001f74
    mem[2014] <= 16'h0613; // 0x80001f78
    mem[2015] <= 16'h2623; // 0x80001f7c
    mem[2016] <= 16'hf0ef; // 0x80001f80
    mem[2017] <= 16'hf06f; // 0x80001f84
    mem[2018] <= 16'h1063; // 0x80001f88
    mem[2019] <= 16'h0493; // 0x80001f8c
    mem[2020] <= 16'hf06f; // 0x80001f90
    mem[2021] <= 16'h1663; // 0x80001f94
    mem[2022] <= 16'h8513; // 0x80001f98
    mem[2023] <= 16'h0593; // 0x80001f9c
    mem[2024] <= 16'hf0ef; // 0x80001fa0
    mem[2025] <= 16'h0593; // 0x80001fa4
    mem[2026] <= 16'h0513; // 0x80001fa8
    mem[2027] <= 16'hf0ef; // 0x80001fac
    mem[2028] <= 16'h0493; // 0x80001fb0
    mem[2029] <= 16'h0593; // 0x80001fb4
    mem[2030] <= 16'hf06f; // 0x80001fb8
    mem[2031] <= 16'h1e63; // 0x80001fbc
    mem[2032] <= 16'h0793; // 0x80001fc0
    mem[2033] <= 16'h2623; // 0x80001fc4
    mem[2034] <= 16'h2c83; // 0x80001fc8
    mem[2035] <= 16'h8063; // 0x80001fcc
    mem[2036] <= 16'h5263; // 0x80001fd0
    mem[2037] <= 16'h0793; // 0x80001fd4
    mem[2038] <= 16'h8463; // 0x80001fd8
    mem[2039] <= 16'h8593; // 0x80001fdc
    mem[2040] <= 16'h8513; // 0x80001fe0
    mem[2041] <= 16'hf0ef; // 0x80001fe4
    mem[2042] <= 16'h0c33; // 0x80001fe8
    mem[2043] <= 16'h5463; // 0x80001fec
    mem[2044] <= 16'h0d13; // 0x80001ff0
    mem[2045] <= 16'h0d13; // 0x80001ff4
    mem[2046] <= 16'h0593; // 0x80001ff8
    mem[2047] <= 16'h8513; // 0x80001ffc
    mem[2048] <= 16'hf0ef; // 0x80002000
    mem[2049] <= 16'h18e3; // 0x80002004
    mem[2050] <= 16'h0793; // 0x80002008
    mem[2051] <= 16'h0c33; // 0x8000200c
    mem[2052] <= 16'h0c33; // 0x80002010
    mem[2053] <= 16'hc503; // 0x80002014
    mem[2054] <= 16'h02e3; // 0x80002018
    mem[2055] <= 16'hc663; // 0x8000201c
    mem[2056] <= 16'h8493; // 0x80002020
    mem[2057] <= 16'h8e63; // 0x80002024
    mem[2058] <= 16'h0593; // 0x80002028
    mem[2059] <= 16'h8c93; // 0x8000202c
    mem[2060] <= 16'hf0ef; // 0x80002030
    mem[2061] <= 16'hc503; // 0x80002034
    mem[2062] <= 16'h0c13; // 0x80002038
    mem[2063] <= 16'h10e3; // 0x8000203c
    mem[2064] <= 16'h5ee3; // 0x80002040
    mem[2065] <= 16'h0493; // 0x80002044
    mem[2066] <= 16'h0c13; // 0x80002048
    mem[2067] <= 16'h0593; // 0x8000204c
    mem[2068] <= 16'h8513; // 0x80002050
    mem[2069] <= 16'hf0ef; // 0x80002054
    mem[2070] <= 16'h18e3; // 0x80002058
    mem[2071] <= 16'hf06f; // 0x8000205c
    mem[2072] <= 16'h1663; // 0x80002060
    mem[2073] <= 16'h0493; // 0x80002064
    mem[2074] <= 16'hf06f; // 0x80002068
    mem[2075] <= 16'h1063; // 0x8000206c
    mem[2076] <= 16'h0513; // 0x80002070
    mem[2077] <= 16'hf0ef; // 0x80002074
    mem[2078] <= 16'h0613; // 0x80002078
    mem[2079] <= 16'h8693; // 0x8000207c
    mem[2080] <= 16'h0493; // 0x80002080
    mem[2081] <= 16'hdce3; // 0x80002084
    mem[2082] <= 16'h2423; // 0x80002088
    mem[2083] <= 16'h2223; // 0x8000208c
    mem[2084] <= 16'h0593; // 0x80002090
    mem[2085] <= 16'h0513; // 0x80002094
    mem[2086] <= 16'hf0ef; // 0x80002098
    mem[2087] <= 16'h2603; // 0x8000209c
    mem[2088] <= 16'h2683; // 0x800020a0
    mem[2089] <= 16'h0633; // 0x800020a4
    mem[2090] <= 16'h37b3; // 0x800020a8
    mem[2091] <= 16'h06b3; // 0x800020ac
    mem[2092] <= 16'h86b3; // 0x800020b0
    mem[2093] <= 16'hf06f; // 0x800020b4
    mem[2094] <= 16'hce03; // 0x800020b8
    mem[2095] <= 16'h8593; // 0x800020bc
    mem[2096] <= 16'h0793; // 0x800020c0
    mem[2097] <= 16'hf06f; // 0x800020c4
    mem[2098] <= 16'h1e63; // 0x800020c8
    mem[2099] <= 16'h0593; // 0x800020cc
    mem[2100] <= 16'h0513; // 0x800020d0
    mem[2101] <= 16'hf0ef; // 0x800020d4
    mem[2102] <= 16'h8413; // 0x800020d8
    mem[2103] <= 16'hf06f; // 0x800020dc
    mem[2104] <= 16'hc503; // 0x800020e0
    mem[2105] <= 16'h1ce3; // 0x800020e4
    mem[2106] <= 16'hf06f; // 0x800020e8
    mem[2107] <= 16'h5463; // 0x800020ec
    mem[2108] <= 16'h0793; // 0x800020f0
    mem[2109] <= 16'h1c97; // 0x800020f4
    mem[2110] <= 16'h8c93; // 0x800020f8
    mem[2111] <= 16'h0513; // 0x800020fc
    mem[2112] <= 16'h9ee3; // 0x80002100
    mem[2113] <= 16'hf06f; // 0x80002104
    mem[2114] <= 16'h8e13; // 0x80002108
    mem[2115] <= 16'h0793; // 0x8000210c
    mem[2116] <= 16'hf06f; // 0x80002110
    mem[2117] <= 16'h0513; // 0x80002114
    mem[2118] <= 16'h1c97; // 0x80002118
    mem[2119] <= 16'h8c93; // 0x8000211c
    mem[2120] <= 16'hf06f; // 0x80002120
    mem[2121] <= 16'h8613; // 0x80002124
    mem[2122] <= 16'hf06f; // 0x80002128
    mem[2123] <= 16'h2623; // 0x8000212c
    mem[2124] <= 16'h0493; // 0x80002130
    mem[2125] <= 16'hf06f; // 0x80002134
    mem[2126] <= 16'h8613; // 0x80002138
    mem[2127] <= 16'hf06f; // 0x8000213c
    mem[2128] <= 16'h2623; // 0x80002140
    mem[2129] <= 16'hf06f; // 0x80002144
    mem[2130] <= 16'h2623; // 0x80002148
    mem[2131] <= 16'h0493; // 0x8000214c
    mem[2132] <= 16'hf06f; // 0x80002150
    mem[2133] <= 16'h2623; // 0x80002154
    mem[2134] <= 16'hf06f; // 0x80002158
    mem[2135] <= 16'h2623; // 0x8000215c
    mem[2136] <= 16'hf06f; // 0x80002160
    mem[2137] <= 16'h2623; // 0x80002164
    mem[2138] <= 16'hf06f; // 0x80002168
    mem[2139] <= 16'h2623; // 0x8000216c
    mem[2140] <= 16'hf06f; // 0x80002170
    mem[2141] <= 16'h0113; // 0x80002174
    mem[2142] <= 16'h0313; // 0x80002178
    mem[2143] <= 16'h2423; // 0x8000217c
    mem[2144] <= 16'h2623; // 0x80002180
    mem[2145] <= 16'h2c23; // 0x80002184
    mem[2146] <= 16'h0413; // 0x80002188
    mem[2147] <= 16'h0613; // 0x8000218c
    mem[2148] <= 16'h0513; // 0x80002190
    mem[2149] <= 16'h2623; // 0x80002194
    mem[2150] <= 16'h2223; // 0x80002198
    mem[2151] <= 16'h2e23; // 0x8000219c
    mem[2152] <= 16'h2023; // 0x800021a0
    mem[2153] <= 16'h2423; // 0x800021a4
    mem[2154] <= 16'h2623; // 0x800021a8
    mem[2155] <= 16'h2e23; // 0x800021ac
    mem[2156] <= 16'hf0ef; // 0x800021b0
    mem[2157] <= 16'h2783; // 0x800021b4
    mem[2158] <= 16'h8023; // 0x800021b8
    mem[2159] <= 16'h2503; // 0x800021bc
    mem[2160] <= 16'h2083; // 0x800021c0
    mem[2161] <= 16'h0533; // 0x800021c4
    mem[2162] <= 16'h2403; // 0x800021c8
    mem[2163] <= 16'h0113; // 0x800021cc
    mem[2164] <= 16'h8067; // 0x800021d0
    mem[2165] <= 16'h0113; // 0x800021d4
    mem[2166] <= 16'h2e23; // 0x800021d8
    mem[2167] <= 16'h2c23; // 0x800021dc
    mem[2168] <= 16'h2a23; // 0x800021e0
    mem[2169] <= 16'h0413; // 0x800021e4
    mem[2170] <= 16'h2823; // 0x800021e8
    mem[2171] <= 16'h2623; // 0x800021ec
    mem[2172] <= 16'h0113; // 0x800021f0
    mem[2173] <= 16'h8993; // 0x800021f4
    mem[2174] <= 16'h0913; // 0x800021f8
    mem[2175] <= 16'hf0ef; // 0x800021fc
    mem[2176] <= 16'h8593; // 0x80002200
    mem[2177] <= 16'h0513; // 0x80002204
    mem[2178] <= 16'hf0ef; // 0x80002208
    mem[2179] <= 16'h0593; // 0x8000220c
    mem[2180] <= 16'h0513; // 0x80002210
    mem[2181] <= 16'h00ef; // 0x80002214
    mem[2182] <= 16'h0493; // 0x80002218
    mem[2183] <= 16'h1697; // 0x8000221c
    mem[2184] <= 16'ha683; // 0x80002220
    mem[2185] <= 16'hf493; // 0x80002224
    mem[2186] <= 16'h0993; // 0x80002228
    mem[2187] <= 16'h9263; // 0x8000222c
    mem[2188] <= 16'h1697; // 0x80002230
    mem[2189] <= 16'ha683; // 0x80002234
    mem[2190] <= 16'h8913; // 0x80002238
    mem[2191] <= 16'h8663; // 0x8000223c
    mem[2192] <= 16'h0513; // 0x80002240
    mem[2193] <= 16'h1617; // 0x80002244
    mem[2194] <= 16'h2603; // 0x80002248
    mem[2195] <= 16'h1597; // 0x8000224c
    mem[2196] <= 16'h8593; // 0x80002250
    mem[2197] <= 16'hf0ef; // 0x80002254
    mem[2198] <= 16'h0933; // 0x80002258
    mem[2199] <= 16'h8663; // 0x8000225c
    mem[2200] <= 16'h8513; // 0x80002260
    mem[2201] <= 16'hf0ef; // 0x80002264
    mem[2202] <= 16'h8513; // 0x80002268
    mem[2203] <= 16'hf0ef; // 0x8000226c
    mem[2204] <= 16'h1617; // 0x80002270
    mem[2205] <= 16'h2603; // 0x80002274
    mem[2206] <= 16'h1597; // 0x80002278
    mem[2207] <= 16'h8593; // 0x8000227c
    mem[2208] <= 16'h8513; // 0x80002280
    mem[2209] <= 16'hf0ef; // 0x80002284
    mem[2210] <= 16'h1697; // 0x80002288
    mem[2211] <= 16'ha683; // 0x8000228c
    mem[2212] <= 16'h8933; // 0x80002290
    mem[2213] <= 16'h84e3; // 0x80002294
    mem[2214] <= 16'hf06f; // 0x80002298
    mem[2215] <= 16'h0113; // 0x8000229c
    mem[2216] <= 16'h2c23; // 0x800022a0
    mem[2217] <= 16'h2823; // 0x800022a4
    mem[2218] <= 16'h2623; // 0x800022a8
    mem[2219] <= 16'h2423; // 0x800022ac
    mem[2220] <= 16'h2223; // 0x800022b0
    mem[2221] <= 16'h2e23; // 0x800022b4
    mem[2222] <= 16'h2a23; // 0x800022b8
    mem[2223] <= 16'h2023; // 0x800022bc
    mem[2224] <= 16'h2e23; // 0x800022c0
    mem[2225] <= 16'h2c23; // 0x800022c4
    mem[2226] <= 16'h2a23; // 0x800022c8
    mem[2227] <= 16'h0413; // 0x800022cc
    mem[2228] <= 16'h2623; // 0x800022d0
    mem[2229] <= 16'h1917; // 0x800022d4
    mem[2230] <= 16'h0913; // 0x800022d8
    mem[2231] <= 16'h0a93; // 0x800022dc
    mem[2232] <= 16'h0a13; // 0x800022e0
    mem[2233] <= 16'h0993; // 0x800022e4
    mem[2234] <= 16'h4503; // 0x800022e8
    mem[2235] <= 16'h0493; // 0x800022ec
    mem[2236] <= 16'h0e63; // 0x800022f0
    mem[2237] <= 16'h0863; // 0x800022f4
    mem[2238] <= 16'h0593; // 0x800022f8
    mem[2239] <= 16'h0413; // 0x800022fc
    mem[2240] <= 16'hf0ef; // 0x80002300
    mem[2241] <= 16'h4503; // 0x80002304
    mem[2242] <= 16'h16e3; // 0x80002308
    mem[2243] <= 16'h2603; // 0x8000230c
    mem[2244] <= 16'h4e03; // 0x80002310
    mem[2245] <= 16'h0c13; // 0x80002314
    mem[2246] <= 16'h0493; // 0x80002318
    mem[2247] <= 16'h0893; // 0x8000231c
    mem[2248] <= 16'h0713; // 0x80002320
    mem[2249] <= 16'h0813; // 0x80002324
    mem[2250] <= 16'h0b13; // 0x80002328
    mem[2251] <= 16'h8b93; // 0x8000232c
    mem[2252] <= 16'h0593; // 0x80002330
    mem[2253] <= 16'h0693; // 0x80002334
    mem[2254] <= 16'h0513; // 0x80002338
    mem[2255] <= 16'h0313; // 0x8000233c
    mem[2256] <= 16'h0793; // 0x80002340
    mem[2257] <= 16'hf793; // 0x80002344
    mem[2258] <= 16'h0413; // 0x80002348
    mem[2259] <= 16'hec63; // 0x8000234c
    mem[2260] <= 16'h9793; // 0x80002350
    mem[2261] <= 16'h87b3; // 0x80002354
    mem[2262] <= 16'ha783; // 0x80002358
    mem[2263] <= 16'h87b3; // 0x8000235c
    mem[2264] <= 16'h8067; // 0x80002360
    mem[2265] <= 16'h2083; // 0x80002364
    mem[2266] <= 16'h2403; // 0x80002368
    mem[2267] <= 16'h2483; // 0x8000236c
    mem[2268] <= 16'h2903; // 0x80002370
    mem[2269] <= 16'h2983; // 0x80002374
    mem[2270] <= 16'h2a03; // 0x80002378
    mem[2271] <= 16'h2a83; // 0x8000237c
    mem[2272] <= 16'h2b03; // 0x80002380
    mem[2273] <= 16'h2b83; // 0x80002384
    mem[2274] <= 16'h2c03; // 0x80002388
    mem[2275] <= 16'h2c83; // 0x8000238c
    mem[2276] <= 16'h0113; // 0x80002390
    mem[2277] <= 16'h8067; // 0x80002394
    mem[2278] <= 16'hd463; // 0x80002398
    mem[2279] <= 16'h0b93; // 0x8000239c
    mem[2280] <= 16'h4e03; // 0x800023a0
    mem[2281] <= 16'h0713; // 0x800023a4
    mem[2282] <= 16'hf06f; // 0x800023a8
    mem[2283] <= 16'h1663; // 0x800023ac
    mem[2284] <= 16'h0c93; // 0x800023b0
    mem[2285] <= 16'h0513; // 0x800023b4
    mem[2286] <= 16'hf0ef; // 0x800023b8
    mem[2287] <= 16'h0c13; // 0x800023bc
    mem[2288] <= 16'h8493; // 0x800023c0
    mem[2289] <= 16'h0713; // 0x800023c4
    mem[2290] <= 16'h8693; // 0x800023c8
    mem[2291] <= 16'h8613; // 0x800023cc
    mem[2292] <= 16'h0513; // 0x800023d0
    mem[2293] <= 16'h8593; // 0x800023d4
    mem[2294] <= 16'hf0ef; // 0x800023d8
    mem[2295] <= 16'hf06f; // 0x800023dc
    mem[2296] <= 16'h1863; // 0x800023e0
    mem[2297] <= 16'h0593; // 0x800023e4
    mem[2298] <= 16'h0513; // 0x800023e8
    mem[2299] <= 16'hf0ef; // 0x800023ec
    mem[2300] <= 16'hf06f; // 0x800023f0
    mem[2301] <= 16'ha483; // 0x800023f4
    mem[2302] <= 16'h4e03; // 0x800023f8
    mem[2303] <= 16'h8893; // 0x800023fc
    mem[2304] <= 16'h0713; // 0x80002400
    mem[2305] <= 16'h8813; // 0x80002404
    mem[2306] <= 16'hdce3; // 0x80002408
    mem[2307] <= 16'h8b93; // 0x8000240c
    mem[2308] <= 16'h0493; // 0x80002410
    mem[2309] <= 16'hf06f; // 0x80002414
    mem[2310] <= 16'h4e03; // 0x80002418
    mem[2311] <= 16'h0b13; // 0x8000241c
    mem[2312] <= 16'h0713; // 0x80002420
    mem[2313] <= 16'hf06f; // 0x80002424
    mem[2314] <= 16'h4e03; // 0x80002428
    mem[2315] <= 16'h0b13; // 0x8000242c
    mem[2316] <= 16'h0713; // 0x80002430
    mem[2317] <= 16'hf06f; // 0x80002434
    mem[2318] <= 16'h4e83; // 0x80002438
    mem[2319] <= 16'h0493; // 0x8000243c
    mem[2320] <= 16'h8793; // 0x80002440
    mem[2321] <= 16'h6063; // 0x80002444
    mem[2322] <= 16'h0713; // 0x80002448
    mem[2323] <= 16'h9793; // 0x8000244c
    mem[2324] <= 16'h84b3; // 0x80002450
    mem[2325] <= 16'h0713; // 0x80002454
    mem[2326] <= 16'h9493; // 0x80002458
    mem[2327] <= 16'h84b3; // 0x8000245c
    mem[2328] <= 16'h4e83; // 0x80002460
    mem[2329] <= 16'h8493; // 0x80002464
    mem[2330] <= 16'h8793; // 0x80002468
    mem[2331] <= 16'h70e3; // 0x8000246c
    mem[2332] <= 16'h8e13; // 0x80002470
    mem[2333] <= 16'hf06f; // 0x80002474
    mem[2334] <= 16'h1463; // 0x80002478
    mem[2335] <= 16'h2503; // 0x8000247c
    mem[2336] <= 16'h0593; // 0x80002480
    mem[2337] <= 16'h0613; // 0x80002484
    mem[2338] <= 16'h2623; // 0x80002488
    mem[2339] <= 16'he0ef; // 0x8000248c
    mem[2340] <= 16'hf06f; // 0x80002490
    mem[2341] <= 16'h1863; // 0x80002494
    mem[2342] <= 16'h0c93; // 0x80002498
    mem[2343] <= 16'hf06f; // 0x8000249c
    mem[2344] <= 16'h1e63; // 0x800024a0
    mem[2345] <= 16'h0593; // 0x800024a4
    mem[2346] <= 16'h0513; // 0x800024a8
    mem[2347] <= 16'he0ef; // 0x800024ac
    mem[2348] <= 16'h0593; // 0x800024b0
    mem[2349] <= 16'h0513; // 0x800024b4
    mem[2350] <= 16'he0ef; // 0x800024b8
    mem[2351] <= 16'h0c93; // 0x800024bc
    mem[2352] <= 16'h0593; // 0x800024c0
    mem[2353] <= 16'hf06f; // 0x800024c4
    mem[2354] <= 16'h1663; // 0x800024c8
    mem[2355] <= 16'h0793; // 0x800024cc
    mem[2356] <= 16'h2623; // 0x800024d0
    mem[2357] <= 16'h2c03; // 0x800024d4
    mem[2358] <= 16'h0863; // 0x800024d8
    mem[2359] <= 16'h5263; // 0x800024dc
    mem[2360] <= 16'h0793; // 0x800024e0
    mem[2361] <= 16'h0c63; // 0x800024e4
    mem[2362] <= 16'h8593; // 0x800024e8
    mem[2363] <= 16'h0513; // 0x800024ec
    mem[2364] <= 16'hf0ef; // 0x800024f0
    mem[2365] <= 16'h8bb3; // 0x800024f4
    mem[2366] <= 16'h5463; // 0x800024f8
    mem[2367] <= 16'h8c93; // 0x800024fc
    mem[2368] <= 16'h8c93; // 0x80002500
    mem[2369] <= 16'h0593; // 0x80002504
    mem[2370] <= 16'h0513; // 0x80002508
    mem[2371] <= 16'he0ef; // 0x8000250c
    mem[2372] <= 16'h98e3; // 0x80002510
    mem[2373] <= 16'h8793; // 0x80002514
    mem[2374] <= 16'h8bb3; // 0x80002518
    mem[2375] <= 16'h8bb3; // 0x8000251c
    mem[2376] <= 16'h4503; // 0x80002520
    mem[2377] <= 16'h02e3; // 0x80002524
    mem[2378] <= 16'hc663; // 0x80002528
    mem[2379] <= 16'h8493; // 0x8000252c
    mem[2380] <= 16'h8e63; // 0x80002530
    mem[2381] <= 16'h0593; // 0x80002534
    mem[2382] <= 16'h0c13; // 0x80002538
    mem[2383] <= 16'he0ef; // 0x8000253c
    mem[2384] <= 16'h4503; // 0x80002540
    mem[2385] <= 16'h8b93; // 0x80002544
    mem[2386] <= 16'h10e3; // 0x80002548
    mem[2387] <= 16'h5ee3; // 0x8000254c
    mem[2388] <= 16'h0493; // 0x80002550
    mem[2389] <= 16'h8b93; // 0x80002554
    mem[2390] <= 16'h0593; // 0x80002558
    mem[2391] <= 16'h8513; // 0x8000255c
    mem[2392] <= 16'he0ef; // 0x80002560
    mem[2393] <= 16'h98e3; // 0x80002564
    mem[2394] <= 16'hf06f; // 0x80002568
    mem[2395] <= 16'h1e63; // 0x8000256c
    mem[2396] <= 16'h0c93; // 0x80002570
    mem[2397] <= 16'hf06f; // 0x80002574
    mem[2398] <= 16'h1863; // 0x80002578
    mem[2399] <= 16'h0513; // 0x8000257c
    mem[2400] <= 16'he0ef; // 0x80002580
    mem[2401] <= 16'h0c13; // 0x80002584
    mem[2402] <= 16'h8493; // 0x80002588
    mem[2403] <= 16'h0c93; // 0x8000258c
    mem[2404] <= 16'hdae3; // 0x80002590
    mem[2405] <= 16'h0593; // 0x80002594
    mem[2406] <= 16'h0513; // 0x80002598
    mem[2407] <= 16'he0ef; // 0x8000259c
    mem[2408] <= 16'h0c33; // 0x800025a0
    mem[2409] <= 16'h37b3; // 0x800025a4
    mem[2410] <= 16'h04b3; // 0x800025a8
    mem[2411] <= 16'h84b3; // 0x800025ac
    mem[2412] <= 16'hf06f; // 0x800025b0
    mem[2413] <= 16'h4e03; // 0x800025b4
    mem[2414] <= 16'h8593; // 0x800025b8
    mem[2415] <= 16'h0713; // 0x800025bc
    mem[2416] <= 16'hf06f; // 0x800025c0
    mem[2417] <= 16'h1e63; // 0x800025c4
    mem[2418] <= 16'h0593; // 0x800025c8
    mem[2419] <= 16'h0513; // 0x800025cc
    mem[2420] <= 16'he0ef; // 0x800025d0
    mem[2421] <= 16'h0413; // 0x800025d4
    mem[2422] <= 16'hf06f; // 0x800025d8
    mem[2423] <= 16'h4503; // 0x800025dc
    mem[2424] <= 16'h14e3; // 0x800025e0
    mem[2425] <= 16'hf06f; // 0x800025e4
    mem[2426] <= 16'h5463; // 0x800025e8
    mem[2427] <= 16'h0793; // 0x800025ec
    mem[2428] <= 16'h1c17; // 0x800025f0
    mem[2429] <= 16'h0c13; // 0x800025f4
    mem[2430] <= 16'h0513; // 0x800025f8
    mem[2431] <= 16'h16e3; // 0x800025fc
    mem[2432] <= 16'hf06f; // 0x80002600
    mem[2433] <= 16'h8e13; // 0x80002604
    mem[2434] <= 16'h0713; // 0x80002608
    mem[2435] <= 16'hf06f; // 0x8000260c
    mem[2436] <= 16'h0513; // 0x80002610
    mem[2437] <= 16'h1c17; // 0x80002614
    mem[2438] <= 16'h0c13; // 0x80002618
    mem[2439] <= 16'hf06f; // 0x8000261c
    mem[2440] <= 16'h8613; // 0x80002620
    mem[2441] <= 16'hf06f; // 0x80002624
    mem[2442] <= 16'h2623; // 0x80002628
    mem[2443] <= 16'h0c93; // 0x8000262c
    mem[2444] <= 16'hf06f; // 0x80002630
    mem[2445] <= 16'h8613; // 0x80002634
    mem[2446] <= 16'hf06f; // 0x80002638
    mem[2447] <= 16'h2623; // 0x8000263c
    mem[2448] <= 16'hf06f; // 0x80002640
    mem[2449] <= 16'h2623; // 0x80002644
    mem[2450] <= 16'h0c93; // 0x80002648
    mem[2451] <= 16'hf06f; // 0x8000264c
    mem[2452] <= 16'h2623; // 0x80002650
    mem[2453] <= 16'hf06f; // 0x80002654
    mem[2454] <= 16'h2623; // 0x80002658
    mem[2455] <= 16'hf06f; // 0x8000265c
    mem[2456] <= 16'h2623; // 0x80002660
    mem[2457] <= 16'hf06f; // 0x80002664
    mem[2458] <= 16'h2623; // 0x80002668
    mem[2459] <= 16'hf06f; // 0x8000266c
    mem[2460] <= 16'h0113; // 0x80002670
    mem[2461] <= 16'h0313; // 0x80002674
    mem[2462] <= 16'h2223; // 0x80002678
    mem[2463] <= 16'h0593; // 0x8000267c
    mem[2464] <= 16'h2e23; // 0x80002680
    mem[2465] <= 16'h2423; // 0x80002684
    mem[2466] <= 16'h2623; // 0x80002688
    mem[2467] <= 16'h2823; // 0x8000268c
    mem[2468] <= 16'h2a23; // 0x80002690
    mem[2469] <= 16'h2c23; // 0x80002694
    mem[2470] <= 16'h2e23; // 0x80002698
    mem[2471] <= 16'h2623; // 0x8000269c
    mem[2472] <= 16'hf0ef; // 0x800026a0
    mem[2473] <= 16'h2083; // 0x800026a4
    mem[2474] <= 16'h0513; // 0x800026a8
    mem[2475] <= 16'h0113; // 0x800026ac
    mem[2476] <= 16'h8067; // 0x800026b0
    mem[2477] <= 16'h0513; // 0x800026b4
    mem[2478] <= 16'h4783; // 0x800026b8
    mem[2479] <= 16'h8593; // 0x800026bc
    mem[2480] <= 16'hc703; // 0x800026c0
    mem[2481] <= 16'h8863; // 0x800026c4
    mem[2482] <= 16'h86e3; // 0x800026c8
    mem[2483] <= 16'h8533; // 0x800026cc
    mem[2484] <= 16'h8067; // 0x800026d0
    mem[2485] <= 16'h0793; // 0x800026d4
    mem[2486] <= 16'hf06f; // 0x800026d8
    mem[2487] <= 16'h0793; // 0x800026dc
    mem[2488] <= 16'h8593; // 0x800026e0
    mem[2489] <= 16'hc703; // 0x800026e4
    mem[2490] <= 16'h8793; // 0x800026e8
    mem[2491] <= 16'h8fa3; // 0x800026ec
    mem[2492] <= 16'h18e3; // 0x800026f0
    mem[2493] <= 16'h8067; // 0x800026f4
    mem[2494] <= 16'h4703; // 0x800026f8
    mem[2495] <= 16'h0693; // 0x800026fc
    mem[2496] <= 16'h0793; // 0x80002700
    mem[2497] <= 16'h1a63; // 0x80002704
    mem[2498] <= 16'h0693; // 0x80002708
    mem[2499] <= 16'h8793; // 0x8000270c
    mem[2500] <= 16'hc703; // 0x80002710
    mem[2501] <= 16'h0ce3; // 0x80002714
    mem[2502] <= 16'h0693; // 0x80002718
    mem[2503] <= 16'hf693; // 0x8000271c
    mem[2504] <= 16'h8063; // 0x80002720
    mem[2505] <= 16'h0593; // 0x80002724
    mem[2506] <= 16'h0a63; // 0x80002728
    mem[2507] <= 16'h0693; // 0x8000272c
    mem[2508] <= 16'h8793; // 0x80002730
    mem[2509] <= 16'h9513; // 0x80002734
    mem[2510] <= 16'h0613; // 0x80002738
    mem[2511] <= 16'hc703; // 0x8000273c
    mem[2512] <= 16'h0533; // 0x80002740
    mem[2513] <= 16'h1513; // 0x80002744
    mem[2514] <= 16'h06b3; // 0x80002748
    mem[2515] <= 16'h12e3; // 0x8000274c
    mem[2516] <= 16'h8463; // 0x80002750
    mem[2517] <= 16'h06b3; // 0x80002754
    mem[2518] <= 16'h8513; // 0x80002758
    mem[2519] <= 16'h8067; // 0x8000275c
    mem[2520] <= 16'h0593; // 0x80002760
    mem[2521] <= 16'hc703; // 0x80002764
    mem[2522] <= 16'hb593; // 0x80002768
    mem[2523] <= 16'h8793; // 0x8000276c
    mem[2524] <= 16'h1ee3; // 0x80002770
    mem[2525] <= 16'h0693; // 0x80002774
    mem[2526] <= 16'hf06f; // 0x80002778
    mem[2527] <= 16'h0693; // 0x8000277c
    mem[2528] <= 16'hf06f; // 0x80002780
    mem[2529] <= 16'h8313; // 0x80002784
    mem[2530] <= 16'h0893; // 0x80002788
    mem[2531] <= 16'h0e13; // 0x8000278c
    mem[2532] <= 16'h8813; // 0x80002790
    mem[2533] <= 16'h9e63; // 0x80002794
    mem[2534] <= 16'hf863; // 0x80002798
    mem[2535] <= 16'h07b7; // 0x8000279c
    mem[2536] <= 16'h7663; // 0x800027a0
    mem[2537] <= 16'h0793; // 0x800027a4
    mem[2538] <= 16'hf463; // 0x800027a8
    mem[2539] <= 16'h0313; // 0x800027ac
    mem[2540] <= 16'h3737; // 0x800027b0
    mem[2541] <= 16'h57b3; // 0x800027b4
    mem[2542] <= 16'h0713; // 0x800027b8
    mem[2543] <= 16'h87b3; // 0x800027bc
    mem[2544] <= 16'hc783; // 0x800027c0
    mem[2545] <= 16'h8333; // 0x800027c4
    mem[2546] <= 16'h0793; // 0x800027c8
    mem[2547] <= 16'h87b3; // 0x800027cc
    mem[2548] <= 16'h8c63; // 0x800027d0
    mem[2549] <= 16'h9733; // 0x800027d4
    mem[2550] <= 16'h5333; // 0x800027d8
    mem[2551] <= 16'h18b3; // 0x800027dc
    mem[2552] <= 16'h6833; // 0x800027e0
    mem[2553] <= 16'h1e33; // 0x800027e4
    mem[2554] <= 16'hd593; // 0x800027e8
    mem[2555] <= 16'h5733; // 0x800027ec
    mem[2556] <= 16'h9613; // 0x800027f0
    mem[2557] <= 16'h5613; // 0x800027f4
    mem[2558] <= 16'h5793; // 0x800027f8
    mem[2559] <= 16'h76b3; // 0x800027fc
    mem[2560] <= 16'h0533; // 0x80002800
    mem[2561] <= 16'h9693; // 0x80002804
    mem[2562] <= 16'he833; // 0x80002808
    mem[2563] <= 16'h7c63; // 0x8000280c
    mem[2564] <= 16'h0833; // 0x80002810
    mem[2565] <= 16'h0793; // 0x80002814
    mem[2566] <= 16'h6463; // 0x80002818
    mem[2567] <= 16'h6863; // 0x8000281c
    mem[2568] <= 16'h8713; // 0x80002820
    mem[2569] <= 16'h0833; // 0x80002824
    mem[2570] <= 16'h5533; // 0x80002828
    mem[2571] <= 16'h1e13; // 0x8000282c
    mem[2572] <= 16'h5e13; // 0x80002830
    mem[2573] <= 16'h7833; // 0x80002834
    mem[2574] <= 16'h0633; // 0x80002838
    mem[2575] <= 16'h1813; // 0x8000283c
    mem[2576] <= 16'h6833; // 0x80002840
    mem[2577] <= 16'h7c63; // 0x80002844
    mem[2578] <= 16'h8833; // 0x80002848
    mem[2579] <= 16'h0793; // 0x8000284c
    mem[2580] <= 16'h6663; // 0x80002850
    mem[2581] <= 16'h0513; // 0x80002854
    mem[2582] <= 16'h7263; // 0x80002858
    mem[2583] <= 16'h1793; // 0x8000285c
    mem[2584] <= 16'he7b3; // 0x80002860
    mem[2585] <= 16'h0593; // 0x80002864
    mem[2586] <= 16'h8513; // 0x80002868
    mem[2587] <= 16'h8067; // 0x8000286c
    mem[2588] <= 16'he663; // 0x80002870
    mem[2589] <= 16'h07b7; // 0x80002874
    mem[2590] <= 16'hea63; // 0x80002878
    mem[2591] <= 16'h0737; // 0x8000287c
    mem[2592] <= 16'h0793; // 0x80002880
    mem[2593] <= 16'hf463; // 0x80002884
    mem[2594] <= 16'h0793; // 0x80002888
    mem[2595] <= 16'h38b7; // 0x8000288c
    mem[2596] <= 16'hd733; // 0x80002890
    mem[2597] <= 16'h8893; // 0x80002894
    mem[2598] <= 16'h0733; // 0x80002898
    mem[2599] <= 16'h4e03; // 0x8000289c
    mem[2600] <= 16'h0e93; // 0x800028a0
    mem[2601] <= 16'h0e33; // 0x800028a4
    mem[2602] <= 16'h8eb3; // 0x800028a8
    mem[2603] <= 16'h9a63; // 0x800028ac
    mem[2604] <= 16'h0593; // 0x800028b0
    mem[2605] <= 16'h0793; // 0x800028b4
    mem[2606] <= 16'h6663; // 0x800028b8
    mem[2607] <= 16'h37b3; // 0x800028bc
    mem[2608] <= 16'hc793; // 0x800028c0
    mem[2609] <= 16'h006f; // 0x800028c4
    mem[2610] <= 16'h1663; // 0x800028c8
    mem[2611] <= 16'h0893; // 0x800028cc
    mem[2612] <= 16'hd8b3; // 0x800028d0
    mem[2613] <= 16'h07b7; // 0x800028d4
    mem[2614] <= 16'he263; // 0x800028d8
    mem[2615] <= 16'h07b7; // 0x800028dc
    mem[2616] <= 16'h0313; // 0x800028e0
    mem[2617] <= 16'hf463; // 0x800028e4
    mem[2618] <= 16'h0313; // 0x800028e8
    mem[2619] <= 16'h3737; // 0x800028ec
    mem[2620] <= 16'hd7b3; // 0x800028f0
    mem[2621] <= 16'h0713; // 0x800028f4
    mem[2622] <= 16'h87b3; // 0x800028f8
    mem[2623] <= 16'hc783; // 0x800028fc
    mem[2624] <= 16'h8333; // 0x80002900
    mem[2625] <= 16'h0793; // 0x80002904
    mem[2626] <= 16'h87b3; // 0x80002908
    mem[2627] <= 16'h9263; // 0x8000290c
    mem[2628] <= 16'h9f13; // 0x80002910
    mem[2629] <= 16'h8733; // 0x80002914
    mem[2630] <= 16'hde93; // 0x80002918
    mem[2631] <= 16'h5f13; // 0x8000291c
    mem[2632] <= 16'h0593; // 0x80002920
    mem[2633] <= 16'h5793; // 0x80002924
    mem[2634] <= 16'h56b3; // 0x80002928
    mem[2635] <= 16'h7733; // 0x8000292c
    mem[2636] <= 16'h8633; // 0x80002930
    mem[2637] <= 16'h1713; // 0x80002934
    mem[2638] <= 16'h67b3; // 0x80002938
    mem[2639] <= 16'hfc63; // 0x8000293c
    mem[2640] <= 16'h87b3; // 0x80002940
    mem[2641] <= 16'h8713; // 0x80002944
    mem[2642] <= 16'he463; // 0x80002948
    mem[2643] <= 16'hea63; // 0x8000294c
    mem[2644] <= 16'h0693; // 0x80002950
    mem[2645] <= 16'h87b3; // 0x80002954
    mem[2646] <= 16'hd533; // 0x80002958
    mem[2647] <= 16'h1e13; // 0x8000295c
    mem[2648] <= 16'h5e13; // 0x80002960
    mem[2649] <= 16'hf7b3; // 0x80002964
    mem[2650] <= 16'h0f33; // 0x80002968
    mem[2651] <= 16'h9793; // 0x8000296c
    mem[2652] <= 16'he7b3; // 0x80002970
    mem[2653] <= 16'hfc63; // 0x80002974
    mem[2654] <= 16'h87b3; // 0x80002978
    mem[2655] <= 16'h0713; // 0x8000297c
    mem[2656] <= 16'hea63; // 0x80002980
    mem[2657] <= 16'h0513; // 0x80002984
    mem[2658] <= 16'hf663; // 0x80002988
    mem[2659] <= 16'h9793; // 0x8000298c
    mem[2660] <= 16'he7b3; // 0x80002990
    mem[2661] <= 16'h8513; // 0x80002994
    mem[2662] <= 16'h8067; // 0x80002998
    mem[2663] <= 16'h0593; // 0x8000299c
    mem[2664] <= 16'h0793; // 0x800029a0
    mem[2665] <= 16'h8513; // 0x800029a4
    mem[2666] <= 16'h8067; // 0x800029a8
    mem[2667] <= 16'h0e13; // 0x800029ac
    mem[2668] <= 16'h37b3; // 0x800029b0
    mem[2669] <= 16'h9793; // 0x800029b4
    mem[2670] <= 16'hf06f; // 0x800029b8
    mem[2671] <= 16'h0793; // 0x800029bc
    mem[2672] <= 16'hf6e3; // 0x800029c0
    mem[2673] <= 16'h0313; // 0x800029c4
    mem[2674] <= 16'hf06f; // 0x800029c8
    mem[2675] <= 16'h07b7; // 0x800029cc
    mem[2676] <= 16'h0313; // 0x800029d0
    mem[2677] <= 16'h7ee3; // 0x800029d4
    mem[2678] <= 16'h0313; // 0x800029d8
    mem[2679] <= 16'hf06f; // 0x800029dc
    mem[2680] <= 16'h5833; // 0x800029e0
    mem[2681] <= 16'h96b3; // 0x800029e4
    mem[2682] <= 16'h6833; // 0x800029e8
    mem[2683] <= 16'hd8b3; // 0x800029ec
    mem[2684] <= 16'h5f13; // 0x800029f0
    mem[2685] <= 16'hd333; // 0x800029f4
    mem[2686] <= 16'h1713; // 0x800029f8
    mem[2687] <= 16'h5713; // 0x800029fc
    mem[2688] <= 16'h95b3; // 0x80002a00
    mem[2689] <= 16'h5e33; // 0x80002a04
    mem[2690] <= 16'h65b3; // 0x80002a08
    mem[2691] <= 16'hd693; // 0x80002a0c
    mem[2692] <= 16'h1633; // 0x80002a10
    mem[2693] <= 16'hf8b3; // 0x80002a14
    mem[2694] <= 16'h07b3; // 0x80002a18
    mem[2695] <= 16'h9893; // 0x80002a1c
    mem[2696] <= 16'he6b3; // 0x80002a20
    mem[2697] <= 16'hfa63; // 0x80002a24
    mem[2698] <= 16'h86b3; // 0x80002a28
    mem[2699] <= 16'h0893; // 0x80002a2c
    mem[2700] <= 16'hf863; // 0x80002a30
    mem[2701] <= 16'h8313; // 0x80002a34
    mem[2702] <= 16'h86b3; // 0x80002a38
    mem[2703] <= 16'hde33; // 0x80002a3c
    mem[2704] <= 16'h9593; // 0x80002a40
    mem[2705] <= 16'hd593; // 0x80002a44
    mem[2706] <= 16'hf6b3; // 0x80002a48
    mem[2707] <= 16'h08b3; // 0x80002a4c
    mem[2708] <= 16'h9693; // 0x80002a50
    mem[2709] <= 16'he733; // 0x80002a54
    mem[2710] <= 16'h7a63; // 0x80002a58
    mem[2711] <= 16'h0733; // 0x80002a5c
    mem[2712] <= 16'h0793; // 0x80002a60
    mem[2713] <= 16'h7663; // 0x80002a64
    mem[2714] <= 16'h8e13; // 0x80002a68
    mem[2715] <= 16'h1793; // 0x80002a6c
    mem[2716] <= 16'h0f37; // 0x80002a70
    mem[2717] <= 16'he7b3; // 0x80002a74
    mem[2718] <= 16'h0693; // 0x80002a78
    mem[2719] <= 16'hf5b3; // 0x80002a7c
    mem[2720] <= 16'hd313; // 0x80002a80
    mem[2721] <= 16'h76b3; // 0x80002a84
    mem[2722] <= 16'h5613; // 0x80002a88
    mem[2723] <= 16'h8e33; // 0x80002a8c
    mem[2724] <= 16'h0733; // 0x80002a90
    mem[2725] <= 16'h85b3; // 0x80002a94
    mem[2726] <= 16'h5813; // 0x80002a98
    mem[2727] <= 16'h06b3; // 0x80002a9c
    mem[2728] <= 16'h85b3; // 0x80002aa0
    mem[2729] <= 16'h05b3; // 0x80002aa4
    mem[2730] <= 16'h0633; // 0x80002aa8
    mem[2731] <= 16'hf463; // 0x80002aac
    mem[2732] <= 16'h0633; // 0x80002ab0
    mem[2733] <= 16'hd693; // 0x80002ab4
    mem[2734] <= 16'h8633; // 0x80002ab8
    mem[2735] <= 16'h6463; // 0x80002abc
    mem[2736] <= 16'h0263; // 0x80002ac0
    mem[2737] <= 16'h0593; // 0x80002ac4
    mem[2738] <= 16'h8513; // 0x80002ac8
    mem[2739] <= 16'h8067; // 0x80002acc
    mem[2740] <= 16'h98b3; // 0x80002ad0
    mem[2741] <= 16'hd633; // 0x80002ad4
    mem[2742] <= 16'hde93; // 0x80002ad8
    mem[2743] <= 16'h5fb3; // 0x80002adc
    mem[2744] <= 16'h9f13; // 0x80002ae0
    mem[2745] <= 16'h5f13; // 0x80002ae4
    mem[2746] <= 16'h9733; // 0x80002ae8
    mem[2747] <= 16'h1e33; // 0x80002aec
    mem[2748] <= 16'h5333; // 0x80002af0
    mem[2749] <= 16'h6733; // 0x80002af4
    mem[2750] <= 16'h5593; // 0x80002af8
    mem[2751] <= 16'h76b3; // 0x80002afc
    mem[2752] <= 16'h07b3; // 0x80002b00
    mem[2753] <= 16'h9693; // 0x80002b04
    mem[2754] <= 16'he6b3; // 0x80002b08
    mem[2755] <= 16'hfe63; // 0x80002b0c
    mem[2756] <= 16'h86b3; // 0x80002b10
    mem[2757] <= 16'h8613; // 0x80002b14
    mem[2758] <= 16'he063; // 0x80002b18
    mem[2759] <= 16'hfe63; // 0x80002b1c
    mem[2760] <= 16'h8f93; // 0x80002b20
    mem[2761] <= 16'h86b3; // 0x80002b24
    mem[2762] <= 16'h86b3; // 0x80002b28
    mem[2763] <= 16'hd7b3; // 0x80002b2c
    mem[2764] <= 16'h1313; // 0x80002b30
    mem[2765] <= 16'h5313; // 0x80002b34
    mem[2766] <= 16'hf6b3; // 0x80002b38
    mem[2767] <= 16'h0633; // 0x80002b3c
    mem[2768] <= 16'h9713; // 0x80002b40
    mem[2769] <= 16'h6733; // 0x80002b44
    mem[2770] <= 16'h7e63; // 0x80002b48
    mem[2771] <= 16'h0733; // 0x80002b4c
    mem[2772] <= 16'h8693; // 0x80002b50
    mem[2773] <= 16'h6e63; // 0x80002b54
    mem[2774] <= 16'h7c63; // 0x80002b58
    mem[2775] <= 16'h8793; // 0x80002b5c
    mem[2776] <= 16'h0733; // 0x80002b60
    mem[2777] <= 16'h9593; // 0x80002b64
    mem[2778] <= 16'h0733; // 0x80002b68
    mem[2779] <= 16'he5b3; // 0x80002b6c
    mem[2780] <= 16'hf06f; // 0x80002b70
    mem[2781] <= 16'h0513; // 0x80002b74
    mem[2782] <= 16'hf06f; // 0x80002b78
    mem[2783] <= 16'h8513; // 0x80002b7c
    mem[2784] <= 16'hf06f; // 0x80002b80
    mem[2785] <= 16'h06b7; // 0x80002b84
    mem[2786] <= 16'h8693; // 0x80002b88
    mem[2787] <= 16'hf733; // 0x80002b8c
    mem[2788] <= 16'h1713; // 0x80002b90
    mem[2789] <= 16'h7e33; // 0x80002b94
    mem[2790] <= 16'h1533; // 0x80002b98
    mem[2791] <= 16'h0733; // 0x80002b9c
    mem[2792] <= 16'h72e3; // 0x80002ba0
    mem[2793] <= 16'h8793; // 0x80002ba4
    mem[2794] <= 16'h0593; // 0x80002ba8
    mem[2795] <= 16'hf06f; // 0x80002bac
    mem[2796] <= 16'h7ce3; // 0x80002bb0
    mem[2797] <= 16'h0e13; // 0x80002bb4
    mem[2798] <= 16'h0733; // 0x80002bb8
    mem[2799] <= 16'hf06f; // 0x80002bbc
    mem[2800] <= 16'hfae3; // 0x80002bc0
    mem[2801] <= 16'h0313; // 0x80002bc4
    mem[2802] <= 16'h86b3; // 0x80002bc8
    mem[2803] <= 16'hf06f; // 0x80002bcc
    mem[2804] <= 16'h8793; // 0x80002bd0
    mem[2805] <= 16'hf06f; // 0x80002bd4
    mem[2806] <= 16'h0f93; // 0x80002bd8
    mem[2807] <= 16'hf06f; // 0x80002bdc
    mem[2808] <= 16'h8693; // 0x80002be0
    mem[2809] <= 16'h87b3; // 0x80002be4
    mem[2810] <= 16'hf06f; // 0x80002be8
    mem[2811] <= 16'h0713; // 0x80002bec
    mem[2812] <= 16'h0833; // 0x80002bf0
    mem[2813] <= 16'hf06f; // 0x80002bf4
    mem[2814] <= 16'h8893; // 0x80002bf8
    mem[2815] <= 16'h0813; // 0x80002bfc
    mem[2816] <= 16'h0e93; // 0x80002c00
    mem[2817] <= 16'h8313; // 0x80002c04
    mem[2818] <= 16'h9863; // 0x80002c08
    mem[2819] <= 16'hfa63; // 0x80002c0c
    mem[2820] <= 16'h07b7; // 0x80002c10
    mem[2821] <= 16'h6c63; // 0x80002c14
    mem[2822] <= 16'h07b7; // 0x80002c18
    mem[2823] <= 16'h0893; // 0x80002c1c
    mem[2824] <= 16'h7463; // 0x80002c20
    mem[2825] <= 16'h0893; // 0x80002c24
    mem[2826] <= 16'h3737; // 0x80002c28
    mem[2827] <= 16'h57b3; // 0x80002c2c
    mem[2828] <= 16'h0713; // 0x80002c30
    mem[2829] <= 16'h87b3; // 0x80002c34
    mem[2830] <= 16'hc783; // 0x80002c38
    mem[2831] <= 16'h0e13; // 0x80002c3c
    mem[2832] <= 16'h88b3; // 0x80002c40
    mem[2833] <= 16'h0e33; // 0x80002c44
    mem[2834] <= 16'h0c63; // 0x80002c48
    mem[2835] <= 16'h95b3; // 0x80002c4c
    mem[2836] <= 16'h58b3; // 0x80002c50
    mem[2837] <= 16'h1833; // 0x80002c54
    mem[2838] <= 16'he333; // 0x80002c58
    mem[2839] <= 16'h1eb3; // 0x80002c5c
    mem[2840] <= 16'h5613; // 0x80002c60
    mem[2841] <= 16'h57b3; // 0x80002c64
    mem[2842] <= 16'h1513; // 0x80002c68
    mem[2843] <= 16'h5513; // 0x80002c6c
    mem[2844] <= 16'hd713; // 0x80002c70
    mem[2845] <= 16'h76b3; // 0x80002c74
    mem[2846] <= 16'h07b3; // 0x80002c78
    mem[2847] <= 16'h9693; // 0x80002c7c
    mem[2848] <= 16'he733; // 0x80002c80
    mem[2849] <= 16'h7863; // 0x80002c84
    mem[2850] <= 16'h0733; // 0x80002c88
    mem[2851] <= 16'h6463; // 0x80002c8c
    mem[2852] <= 16'h6c63; // 0x80002c90
    mem[2853] <= 16'h0733; // 0x80002c94
    mem[2854] <= 16'h56b3; // 0x80002c98
    mem[2855] <= 16'h9793; // 0x80002c9c
    mem[2856] <= 16'hd793; // 0x80002ca0
    mem[2857] <= 16'h7733; // 0x80002ca4
    mem[2858] <= 16'h0533; // 0x80002ca8
    mem[2859] <= 16'h1713; // 0x80002cac
    mem[2860] <= 16'h67b3; // 0x80002cb0
    mem[2861] <= 16'hfa63; // 0x80002cb4
    mem[2862] <= 16'h87b3; // 0x80002cb8
    mem[2863] <= 16'he663; // 0x80002cbc
    mem[2864] <= 16'hf463; // 0x80002cc0
    mem[2865] <= 16'h87b3; // 0x80002cc4
    mem[2866] <= 16'h8533; // 0x80002cc8
    mem[2867] <= 16'h5533; // 0x80002ccc
    mem[2868] <= 16'h0593; // 0x80002cd0
    mem[2869] <= 16'h8067; // 0x80002cd4
    mem[2870] <= 16'heee3; // 0x80002cd8
    mem[2871] <= 16'h07b7; // 0x80002cdc
    mem[2872] <= 16'he663; // 0x80002ce0
    mem[2873] <= 16'h0737; // 0x80002ce4
    mem[2874] <= 16'h0793; // 0x80002ce8
    mem[2875] <= 16'hf463; // 0x80002cec
    mem[2876] <= 16'h0793; // 0x80002cf0
    mem[2877] <= 16'h3e37; // 0x80002cf4
    mem[2878] <= 16'h0e13; // 0x80002cf8
    mem[2879] <= 16'hd733; // 0x80002cfc
    mem[2880] <= 16'h0733; // 0x80002d00
    mem[2881] <= 16'h4f03; // 0x80002d04
    mem[2882] <= 16'h0e13; // 0x80002d08
    mem[2883] <= 16'h0f33; // 0x80002d0c
    mem[2884] <= 16'h0e33; // 0x80002d10
    mem[2885] <= 16'h1463; // 0x80002d14
    mem[2886] <= 16'he663; // 0x80002d18
    mem[2887] <= 16'h0793; // 0x80002d1c
    mem[2888] <= 16'hea63; // 0x80002d20
    mem[2889] <= 16'h07b3; // 0x80002d24
    mem[2890] <= 16'h85b3; // 0x80002d28
    mem[2891] <= 16'h36b3; // 0x80002d2c
    mem[2892] <= 16'h8333; // 0x80002d30
    mem[2893] <= 16'h8513; // 0x80002d34
    mem[2894] <= 16'h0593; // 0x80002d38
    mem[2895] <= 16'h8067; // 0x80002d3c
    mem[2896] <= 16'h1663; // 0x80002d40
    mem[2897] <= 16'h0813; // 0x80002d44
    mem[2898] <= 16'h5833; // 0x80002d48
    mem[2899] <= 16'h07b7; // 0x80002d4c
    mem[2900] <= 16'h6663; // 0x80002d50
    mem[2901] <= 16'h07b7; // 0x80002d54
    mem[2902] <= 16'h0893; // 0x80002d58
    mem[2903] <= 16'h7463; // 0x80002d5c
    mem[2904] <= 16'h0893; // 0x80002d60
    mem[2905] <= 16'h3737; // 0x80002d64
    mem[2906] <= 16'h57b3; // 0x80002d68
    mem[2907] <= 16'h0713; // 0x80002d6c
    mem[2908] <= 16'h87b3; // 0x80002d70
    mem[2909] <= 16'hc783; // 0x80002d74
    mem[2910] <= 16'h0e13; // 0x80002d78
    mem[2911] <= 16'h88b3; // 0x80002d7c
    mem[2912] <= 16'h0e33; // 0x80002d80
    mem[2913] <= 16'h1063; // 0x80002d84
    mem[2914] <= 16'h1793; // 0x80002d88
    mem[2915] <= 16'h85b3; // 0x80002d8c
    mem[2916] <= 16'h5613; // 0x80002d90
    mem[2917] <= 16'hd793; // 0x80002d94
    mem[2918] <= 16'hd713; // 0x80002d98
    mem[2919] <= 16'hd6b3; // 0x80002d9c
    mem[2920] <= 16'hf5b3; // 0x80002da0
    mem[2921] <= 16'h86b3; // 0x80002da4
    mem[2922] <= 16'h9593; // 0x80002da8
    mem[2923] <= 16'he733; // 0x80002dac
    mem[2924] <= 16'h7a63; // 0x80002db0
    mem[2925] <= 16'h0733; // 0x80002db4
    mem[2926] <= 16'h6663; // 0x80002db8
    mem[2927] <= 16'h7463; // 0x80002dbc
    mem[2928] <= 16'h0733; // 0x80002dc0
    mem[2929] <= 16'h0733; // 0x80002dc4
    mem[2930] <= 16'h5533; // 0x80002dc8
    mem[2931] <= 16'h9e93; // 0x80002dcc
    mem[2932] <= 16'hde93; // 0x80002dd0
    mem[2933] <= 16'h7733; // 0x80002dd4
    mem[2934] <= 16'h0533; // 0x80002dd8
    mem[2935] <= 16'h1713; // 0x80002ddc
    mem[2936] <= 16'h67b3; // 0x80002de0
    mem[2937] <= 16'hf2e3; // 0x80002de4
    mem[2938] <= 16'hf06f; // 0x80002de8
    mem[2939] <= 16'h0f13; // 0x80002dec
    mem[2940] <= 16'h37b3; // 0x80002df0
    mem[2941] <= 16'h9793; // 0x80002df4
    mem[2942] <= 16'hf06f; // 0x80002df8
    mem[2943] <= 16'h0793; // 0x80002dfc
    mem[2944] <= 16'hf2e3; // 0x80002e00
    mem[2945] <= 16'h0893; // 0x80002e04
    mem[2946] <= 16'hf06f; // 0x80002e08
    mem[2947] <= 16'h0793; // 0x80002e0c
    mem[2948] <= 16'hfce3; // 0x80002e10
    mem[2949] <= 16'h0893; // 0x80002e14
    mem[2950] <= 16'hf06f; // 0x80002e18
    mem[2951] <= 16'h57b3; // 0x80002e1c
    mem[2952] <= 16'h96b3; // 0x80002e20
    mem[2953] <= 16'he6b3; // 0x80002e24
    mem[2954] <= 16'hd8b3; // 0x80002e28
    mem[2955] <= 16'hd713; // 0x80002e2c
    mem[2956] <= 16'hd333; // 0x80002e30
    mem[2957] <= 16'h9f93; // 0x80002e34
    mem[2958] <= 16'h57b3; // 0x80002e38
    mem[2959] <= 16'hdf93; // 0x80002e3c
    mem[2960] <= 16'h95b3; // 0x80002e40
    mem[2961] <= 16'he5b3; // 0x80002e44
    mem[2962] <= 16'h17b3; // 0x80002e48
    mem[2963] <= 16'hd813; // 0x80002e4c
    mem[2964] <= 16'h1533; // 0x80002e50
    mem[2965] <= 16'hf8b3; // 0x80002e54
    mem[2966] <= 16'h8633; // 0x80002e58
    mem[2967] <= 16'h9893; // 0x80002e5c
    mem[2968] <= 16'he833; // 0x80002e60
    mem[2969] <= 16'h7a63; // 0x80002e64
    mem[2970] <= 16'h0833; // 0x80002e68
    mem[2971] <= 16'h0893; // 0x80002e6c
    mem[2972] <= 16'h7463; // 0x80002e70
    mem[2973] <= 16'h8313; // 0x80002e74
    mem[2974] <= 16'h0833; // 0x80002e78
    mem[2975] <= 16'h5633; // 0x80002e7c
    mem[2976] <= 16'h9593; // 0x80002e80
    mem[2977] <= 16'hd593; // 0x80002e84
    mem[2978] <= 16'h7833; // 0x80002e88
    mem[2979] <= 16'h8fb3; // 0x80002e8c
    mem[2980] <= 16'h1713; // 0x80002e90
    mem[2981] <= 16'h6733; // 0x80002e94
    mem[2982] <= 16'h7a63; // 0x80002e98
    mem[2983] <= 16'h0733; // 0x80002e9c
    mem[2984] <= 16'h0593; // 0x80002ea0
    mem[2985] <= 16'h7263; // 0x80002ea4
    mem[2986] <= 16'h8613; // 0x80002ea8
    mem[2987] <= 16'h1313; // 0x80002eac
    mem[2988] <= 16'h05b7; // 0x80002eb0
    mem[2989] <= 16'h6333; // 0x80002eb4
    mem[2990] <= 16'h8893; // 0x80002eb8
    mem[2991] <= 16'h7eb3; // 0x80002ebc
    mem[2992] <= 16'hd613; // 0x80002ec0
    mem[2993] <= 16'h5313; // 0x80002ec4
    mem[2994] <= 16'hf8b3; // 0x80002ec8
    mem[2995] <= 16'h82b3; // 0x80002ecc
    mem[2996] <= 16'h0733; // 0x80002ed0
    mem[2997] <= 16'h8eb3; // 0x80002ed4
    mem[2998] <= 16'hd813; // 0x80002ed8
    mem[2999] <= 16'h08b3; // 0x80002edc
    mem[3000] <= 16'h8eb3; // 0x80002ee0
    mem[3001] <= 16'h0833; // 0x80002ee4
    mem[3002] <= 16'h0633; // 0x80002ee8
    mem[3003] <= 16'h7463; // 0x80002eec
    mem[3004] <= 16'h0633; // 0x80002ef0
    mem[3005] <= 16'h08b7; // 0x80002ef4
    mem[3006] <= 16'h8893; // 0x80002ef8
    mem[3007] <= 16'h5593; // 0x80002efc
    mem[3008] <= 16'h7833; // 0x80002f00
    mem[3009] <= 16'h1813; // 0x80002f04
    mem[3010] <= 16'hf2b3; // 0x80002f08
    mem[3011] <= 16'h8633; // 0x80002f0c
    mem[3012] <= 16'h0833; // 0x80002f10
    mem[3013] <= 16'h6e63; // 0x80002f14
    mem[3014] <= 16'h0c63; // 0x80002f18
    mem[3015] <= 16'h05b3; // 0x80002f1c
    mem[3016] <= 16'h0793; // 0x80002f20
    mem[3017] <= 16'h07b3; // 0x80002f24
    mem[3018] <= 16'h3533; // 0x80002f28
    mem[3019] <= 16'h85b3; // 0x80002f2c
    mem[3020] <= 16'h9f33; // 0x80002f30
    mem[3021] <= 16'hd533; // 0x80002f34
    mem[3022] <= 16'h6533; // 0x80002f38
    mem[3023] <= 16'hd5b3; // 0x80002f3c
    mem[3024] <= 16'h8067; // 0x80002f40
    mem[3025] <= 16'h1833; // 0x80002f44
    mem[3026] <= 16'hd733; // 0x80002f48
    mem[3027] <= 16'h5613; // 0x80002f4c
    mem[3028] <= 16'h56b3; // 0x80002f50
    mem[3029] <= 16'h1793; // 0x80002f54
    mem[3030] <= 16'hd793; // 0x80002f58
    mem[3031] <= 16'h58b3; // 0x80002f5c
    mem[3032] <= 16'h1eb3; // 0x80002f60
    mem[3033] <= 16'h95b3; // 0x80002f64
    mem[3034] <= 16'he5b3; // 0x80002f68
    mem[3035] <= 16'hd893; // 0x80002f6c
    mem[3036] <= 16'h7733; // 0x80002f70
    mem[3037] <= 16'h8533; // 0x80002f74
    mem[3038] <= 16'h1693; // 0x80002f78
    mem[3039] <= 16'he6b3; // 0x80002f7c
    mem[3040] <= 16'hfa63; // 0x80002f80
    mem[3041] <= 16'h86b3; // 0x80002f84
    mem[3042] <= 16'he663; // 0x80002f88
    mem[3043] <= 16'hf463; // 0x80002f8c
    mem[3044] <= 16'h86b3; // 0x80002f90
    mem[3045] <= 16'h86b3; // 0x80002f94
    mem[3046] <= 16'hd733; // 0x80002f98
    mem[3047] <= 16'h9893; // 0x80002f9c
    mem[3048] <= 16'hd893; // 0x80002fa0
    mem[3049] <= 16'hf6b3; // 0x80002fa4
    mem[3050] <= 16'h8733; // 0x80002fa8
    mem[3051] <= 16'h9593; // 0x80002fac
    mem[3052] <= 16'he5b3; // 0x80002fb0
    mem[3053] <= 16'hfa63; // 0x80002fb4
    mem[3054] <= 16'h85b3; // 0x80002fb8
    mem[3055] <= 16'he663; // 0x80002fbc
    mem[3056] <= 16'hf463; // 0x80002fc0
    mem[3057] <= 16'h85b3; // 0x80002fc4
    mem[3058] <= 16'h85b3; // 0x80002fc8
    mem[3059] <= 16'hf06f; // 0x80002fcc
    mem[3060] <= 16'h07b3; // 0x80002fd0
    mem[3061] <= 16'h05b3; // 0x80002fd4
    mem[3062] <= 16'h3833; // 0x80002fd8
    mem[3063] <= 16'h85b3; // 0x80002fdc
    mem[3064] <= 16'h05b3; // 0x80002fe0
    mem[3065] <= 16'hf06f; // 0x80002fe4
    mem[3066] <= 16'h70e3; // 0x80002fe8
    mem[3067] <= 16'h0613; // 0x80002fec
    mem[3068] <= 16'h0733; // 0x80002ff0
    mem[3069] <= 16'hf06f; // 0x80002ff4
    mem[3070] <= 16'h7ee3; // 0x80002ff8
    mem[3071] <= 16'h0313; // 0x80002ffc
    mem[3072] <= 16'h0833; // 0x80003000
    mem[3073] <= 16'hf06f; // 0x80003004
    mem[3074] <= 16'h0733; // 0x80003008
    mem[3075] <= 16'hf06f; // 0x8000300c
    mem[3076] <= 16'h60e3; // 0x80003010
    mem[3077] <= 16'h0793; // 0x80003014
    mem[3078] <= 16'h0593; // 0x80003018
    mem[3079] <= 16'hf06f; // 0x8000301c
    mem[3080] <= 16'h0613; // 0x80003020
    mem[3081] <= 16'h0513; // 0x80003024
    mem[3082] <= 16'hf693; // 0x80003028
    mem[3083] <= 16'h8463; // 0x8000302c
    mem[3084] <= 16'h0533; // 0x80003030
    mem[3085] <= 16'hd593; // 0x80003034
    mem[3086] <= 16'h1613; // 0x80003038
    mem[3087] <= 16'h96e3; // 0x8000303c
    mem[3088] <= 16'h8067; // 0x80003040
 
 
//================================================================
//== Section  .text.startup
//================================================================
    mem[3089] <= 16'h07b7; // 0x80003044
    mem[3090] <= 16'h0713; // 0x80003048
    mem[3091] <= 16'ha683; // 0x8000304c
    mem[3092] <= 16'h5ee3; // 0x80003050
    mem[3093] <= 16'h0713; // 0x80003054
    mem[3094] <= 16'ha423; // 0x80003058
    mem[3095] <= 16'h0793; // 0x8000305c
    mem[3096] <= 16'ha7f3; // 0x80003060
    mem[3097] <= 16'h006f; // 0x80003064
    mem[3098] <= 16'h0113; // 0x80003068
    mem[3099] <= 16'h0517; // 0x8000306c
    mem[3100] <= 16'h0513; // 0x80003070
    mem[3101] <= 16'h2623; // 0x80003074
    mem[3102] <= 16'hf317; // 0x80003078
    mem[3103] <= 16'h00e7; // 0x8000307c
    mem[3104] <= 16'h2083; // 0x80003080
    mem[3105] <= 16'h0513; // 0x80003084
    mem[3106] <= 16'h0113; // 0x80003088
    mem[3107] <= 16'h8067; // 0x8000308c
 
 
//================================================================
//== Section  .rodata
//================================================================
    mem[3108] <= 16'hee08; // 0x80003090
    mem[3109] <= 16'hf038; // 0x80003094
    mem[3110] <= 16'hee44; // 0x80003098
    mem[3111] <= 16'hf038; // 0x8000309c
    mem[3112] <= 16'hf038; // 0x800030a0
    mem[3113] <= 16'hf038; // 0x800030a4
    mem[3114] <= 16'hf038; // 0x800030a8
    mem[3115] <= 16'hee58; // 0x800030ac
    mem[3116] <= 16'hf038; // 0x800030b0
    mem[3117] <= 16'hf038; // 0x800030b4
    mem[3118] <= 16'hee7c; // 0x800030b8
    mem[3119] <= 16'hee00; // 0x800030bc
    mem[3120] <= 16'hf038; // 0x800030c0
    mem[3121] <= 16'hee8c; // 0x800030c4
    mem[3122] <= 16'hee9c; // 0x800030c8
    mem[3123] <= 16'hee9c; // 0x800030cc
    mem[3124] <= 16'hee9c; // 0x800030d0
    mem[3125] <= 16'hee9c; // 0x800030d4
    mem[3126] <= 16'hee9c; // 0x800030d8
    mem[3127] <= 16'hee9c; // 0x800030dc
    mem[3128] <= 16'hee9c; // 0x800030e0
    mem[3129] <= 16'hee9c; // 0x800030e4
    mem[3130] <= 16'hee9c; // 0x800030e8
    mem[3131] <= 16'hf038; // 0x800030ec
    mem[3132] <= 16'hf038; // 0x800030f0
    mem[3133] <= 16'hf038; // 0x800030f4
    mem[3134] <= 16'hf038; // 0x800030f8
    mem[3135] <= 16'hf038; // 0x800030fc
    mem[3136] <= 16'hf038; // 0x80003100
    mem[3137] <= 16'hf038; // 0x80003104
    mem[3138] <= 16'hf038; // 0x80003108
    mem[3139] <= 16'hf038; // 0x8000310c
    mem[3140] <= 16'hf038; // 0x80003110
    mem[3141] <= 16'hf038; // 0x80003114
    mem[3142] <= 16'hf038; // 0x80003118
    mem[3143] <= 16'hf038; // 0x8000311c
    mem[3144] <= 16'hf038; // 0x80003120
    mem[3145] <= 16'hf038; // 0x80003124
    mem[3146] <= 16'hf038; // 0x80003128
    mem[3147] <= 16'hf038; // 0x8000312c
    mem[3148] <= 16'hf038; // 0x80003130
    mem[3149] <= 16'hf038; // 0x80003134
    mem[3150] <= 16'hf038; // 0x80003138
    mem[3151] <= 16'hf038; // 0x8000313c
    mem[3152] <= 16'hf038; // 0x80003140
    mem[3153] <= 16'hf038; // 0x80003144
    mem[3154] <= 16'hf038; // 0x80003148
    mem[3155] <= 16'hf038; // 0x8000314c
    mem[3156] <= 16'hf038; // 0x80003150
    mem[3157] <= 16'hf038; // 0x80003154
    mem[3158] <= 16'hf038; // 0x80003158
    mem[3159] <= 16'hf038; // 0x8000315c
    mem[3160] <= 16'hf038; // 0x80003160
    mem[3161] <= 16'hf038; // 0x80003164
    mem[3162] <= 16'hf038; // 0x80003168
    mem[3163] <= 16'hf038; // 0x8000316c
    mem[3164] <= 16'hf038; // 0x80003170
    mem[3165] <= 16'hf038; // 0x80003174
    mem[3166] <= 16'hf038; // 0x80003178
    mem[3167] <= 16'hf038; // 0x8000317c
    mem[3168] <= 16'hf038; // 0x80003180
    mem[3169] <= 16'hf038; // 0x80003184
    mem[3170] <= 16'hf038; // 0x80003188
    mem[3171] <= 16'hf038; // 0x8000318c
    mem[3172] <= 16'heedc; // 0x80003190
    mem[3173] <= 16'hefdc; // 0x80003194
    mem[3174] <= 16'hf038; // 0x80003198
    mem[3175] <= 16'hf038; // 0x8000319c
    mem[3176] <= 16'hf038; // 0x800031a0
    mem[3177] <= 16'hf038; // 0x800031a4
    mem[3178] <= 16'hf038; // 0x800031a8
    mem[3179] <= 16'hf038; // 0x800031ac
    mem[3180] <= 16'hf038; // 0x800031b0
    mem[3181] <= 16'hf028; // 0x800031b4
    mem[3182] <= 16'hf038; // 0x800031b8
    mem[3183] <= 16'hf038; // 0x800031bc
    mem[3184] <= 16'heef8; // 0x800031c0
    mem[3185] <= 16'hef04; // 0x800031c4
    mem[3186] <= 16'hf038; // 0x800031c8
    mem[3187] <= 16'hf038; // 0x800031cc
    mem[3188] <= 16'hef2c; // 0x800031d0
    mem[3189] <= 16'hf038; // 0x800031d4
    mem[3190] <= 16'hefd0; // 0x800031d8
    mem[3191] <= 16'hf038; // 0x800031dc
    mem[3192] <= 16'hf038; // 0x800031e0
    mem[3193] <= 16'hee14; // 0x800031e4
    mem[3194] <= 16'hf1b8; // 0x800031e8
    mem[3195] <= 16'hf3dc; // 0x800031ec
    mem[3196] <= 16'hf1f8; // 0x800031f0
    mem[3197] <= 16'hf3dc; // 0x800031f4
    mem[3198] <= 16'hf3dc; // 0x800031f8
    mem[3199] <= 16'hf3dc; // 0x800031fc
    mem[3200] <= 16'hf3dc; // 0x80003200
    mem[3201] <= 16'hf20c; // 0x80003204
    mem[3202] <= 16'hf3dc; // 0x80003208
    mem[3203] <= 16'hf3dc; // 0x8000320c
    mem[3204] <= 16'hf230; // 0x80003210
    mem[3205] <= 16'hf1b0; // 0x80003214
    mem[3206] <= 16'hf3dc; // 0x80003218
    mem[3207] <= 16'hf240; // 0x8000321c
    mem[3208] <= 16'hf250; // 0x80003220
    mem[3209] <= 16'hf250; // 0x80003224
    mem[3210] <= 16'hf250; // 0x80003228
    mem[3211] <= 16'hf250; // 0x8000322c
    mem[3212] <= 16'hf250; // 0x80003230
    mem[3213] <= 16'hf250; // 0x80003234
    mem[3214] <= 16'hf250; // 0x80003238
    mem[3215] <= 16'hf250; // 0x8000323c
    mem[3216] <= 16'hf250; // 0x80003240
    mem[3217] <= 16'hf3dc; // 0x80003244
    mem[3218] <= 16'hf3dc; // 0x80003248
    mem[3219] <= 16'hf3dc; // 0x8000324c
    mem[3220] <= 16'hf3dc; // 0x80003250
    mem[3221] <= 16'hf3dc; // 0x80003254
    mem[3222] <= 16'hf3dc; // 0x80003258
    mem[3223] <= 16'hf3dc; // 0x8000325c
    mem[3224] <= 16'hf3dc; // 0x80003260
    mem[3225] <= 16'hf3dc; // 0x80003264
    mem[3226] <= 16'hf3dc; // 0x80003268
    mem[3227] <= 16'hf3dc; // 0x8000326c
    mem[3228] <= 16'hf3dc; // 0x80003270
    mem[3229] <= 16'hf3dc; // 0x80003274
    mem[3230] <= 16'hf3dc; // 0x80003278
    mem[3231] <= 16'hf3dc; // 0x8000327c
    mem[3232] <= 16'hf3dc; // 0x80003280
    mem[3233] <= 16'hf3dc; // 0x80003284
    mem[3234] <= 16'hf3dc; // 0x80003288
    mem[3235] <= 16'hf3dc; // 0x8000328c
    mem[3236] <= 16'hf3dc; // 0x80003290
    mem[3237] <= 16'hf3dc; // 0x80003294
    mem[3238] <= 16'hf3dc; // 0x80003298
    mem[3239] <= 16'hf3dc; // 0x8000329c
    mem[3240] <= 16'hf3dc; // 0x800032a0
    mem[3241] <= 16'hf3dc; // 0x800032a4
    mem[3242] <= 16'hf3dc; // 0x800032a8
    mem[3243] <= 16'hf3dc; // 0x800032ac
    mem[3244] <= 16'hf3dc; // 0x800032b0
    mem[3245] <= 16'hf3dc; // 0x800032b4
    mem[3246] <= 16'hf3dc; // 0x800032b8
    mem[3247] <= 16'hf3dc; // 0x800032bc
    mem[3248] <= 16'hf3dc; // 0x800032c0
    mem[3249] <= 16'hf3dc; // 0x800032c4
    mem[3250] <= 16'hf3dc; // 0x800032c8
    mem[3251] <= 16'hf3dc; // 0x800032cc
    mem[3252] <= 16'hf3dc; // 0x800032d0
    mem[3253] <= 16'hf3dc; // 0x800032d4
    mem[3254] <= 16'hf3dc; // 0x800032d8
    mem[3255] <= 16'hf3dc; // 0x800032dc
    mem[3256] <= 16'hf3dc; // 0x800032e0
    mem[3257] <= 16'hf3dc; // 0x800032e4
    mem[3258] <= 16'hf290; // 0x800032e8
    mem[3259] <= 16'hf390; // 0x800032ec
    mem[3260] <= 16'hf3dc; // 0x800032f0
    mem[3261] <= 16'hf3dc; // 0x800032f4
    mem[3262] <= 16'hf3dc; // 0x800032f8
    mem[3263] <= 16'hf3dc; // 0x800032fc
    mem[3264] <= 16'hf3dc; // 0x80003300
    mem[3265] <= 16'hf3dc; // 0x80003304
    mem[3266] <= 16'hf3dc; // 0x80003308
    mem[3267] <= 16'hf3cc; // 0x8000330c
    mem[3268] <= 16'hf3dc; // 0x80003310
    mem[3269] <= 16'hf3dc; // 0x80003314
    mem[3270] <= 16'hf2ac; // 0x80003318
    mem[3271] <= 16'hf2b8; // 0x8000331c
    mem[3272] <= 16'hf3dc; // 0x80003320
    mem[3273] <= 16'hf3dc; // 0x80003324
    mem[3274] <= 16'hf2e0; // 0x80003328
    mem[3275] <= 16'hf3dc; // 0x8000332c
    mem[3276] <= 16'hf384; // 0x80003330
    mem[3277] <= 16'hf3dc; // 0x80003334
    mem[3278] <= 16'hf3dc; // 0x80003338
    mem[3279] <= 16'hf1c4; // 0x8000333c
    mem[3280] <= 16'h0100; // 0x80003340
    mem[3281] <= 16'h0303; // 0x80003344
    mem[3282] <= 16'h0404; // 0x80003348
    mem[3283] <= 16'h0404; // 0x8000334c
    mem[3284] <= 16'h0505; // 0x80003350
    mem[3285] <= 16'h0505; // 0x80003354
    mem[3286] <= 16'h0505; // 0x80003358
    mem[3287] <= 16'h0505; // 0x8000335c
    mem[3288] <= 16'h0606; // 0x80003360
    mem[3289] <= 16'h0606; // 0x80003364
    mem[3290] <= 16'h0606; // 0x80003368
    mem[3291] <= 16'h0606; // 0x8000336c
    mem[3292] <= 16'h0606; // 0x80003370
    mem[3293] <= 16'h0606; // 0x80003374
    mem[3294] <= 16'h0606; // 0x80003378
    mem[3295] <= 16'h0606; // 0x8000337c
    mem[3296] <= 16'h0707; // 0x80003380
    mem[3297] <= 16'h0707; // 0x80003384
    mem[3298] <= 16'h0707; // 0x80003388
    mem[3299] <= 16'h0707; // 0x8000338c
    mem[3300] <= 16'h0707; // 0x80003390
    mem[3301] <= 16'h0707; // 0x80003394
    mem[3302] <= 16'h0707; // 0x80003398
    mem[3303] <= 16'h0707; // 0x8000339c
    mem[3304] <= 16'h0707; // 0x800033a0
    mem[3305] <= 16'h0707; // 0x800033a4
    mem[3306] <= 16'h0707; // 0x800033a8
    mem[3307] <= 16'h0707; // 0x800033ac
    mem[3308] <= 16'h0707; // 0x800033b0
    mem[3309] <= 16'h0707; // 0x800033b4
    mem[3310] <= 16'h0707; // 0x800033b8
    mem[3311] <= 16'h0707; // 0x800033bc
    mem[3312] <= 16'h0808; // 0x800033c0
    mem[3313] <= 16'h0808; // 0x800033c4
    mem[3314] <= 16'h0808; // 0x800033c8
    mem[3315] <= 16'h0808; // 0x800033cc
    mem[3316] <= 16'h0808; // 0x800033d0
    mem[3317] <= 16'h0808; // 0x800033d4
    mem[3318] <= 16'h0808; // 0x800033d8
    mem[3319] <= 16'h0808; // 0x800033dc
    mem[3320] <= 16'h0808; // 0x800033e0
    mem[3321] <= 16'h0808; // 0x800033e4
    mem[3322] <= 16'h0808; // 0x800033e8
    mem[3323] <= 16'h0808; // 0x800033ec
    mem[3324] <= 16'h0808; // 0x800033f0
    mem[3325] <= 16'h0808; // 0x800033f4
    mem[3326] <= 16'h0808; // 0x800033f8
    mem[3327] <= 16'h0808; // 0x800033fc
    mem[3328] <= 16'h0808; // 0x80003400
    mem[3329] <= 16'h0808; // 0x80003404
    mem[3330] <= 16'h0808; // 0x80003408
    mem[3331] <= 16'h0808; // 0x8000340c
    mem[3332] <= 16'h0808; // 0x80003410
    mem[3333] <= 16'h0808; // 0x80003414
    mem[3334] <= 16'h0808; // 0x80003418
    mem[3335] <= 16'h0808; // 0x8000341c
    mem[3336] <= 16'h0808; // 0x80003420
    mem[3337] <= 16'h0808; // 0x80003424
    mem[3338] <= 16'h0808; // 0x80003428
    mem[3339] <= 16'h0808; // 0x8000342c
    mem[3340] <= 16'h0808; // 0x80003430
    mem[3341] <= 16'h0808; // 0x80003434
    mem[3342] <= 16'h0808; // 0x80003438
    mem[3343] <= 16'h0808; // 0x8000343c
 
 
//================================================================
//== Section  .rodata.str1.4
//================================================================
    mem[3344] <= 16'h636d; // 0x80003440
    mem[3345] <= 16'h656c; // 0x80003444
    mem[3346] <= 16'h696d; // 0x80003448
    mem[3347] <= 16'h7274; // 0x8000344c
    mem[3348] <= 16'h0000; // 0x80003450
    mem[3349] <= 16'h6d49; // 0x80003454
    mem[3350] <= 16'h6d65; // 0x80003458
    mem[3351] <= 16'h2074; // 0x8000345c
    mem[3352] <= 16'h6e69; // 0x80003460
    mem[3353] <= 16'h202c; // 0x80003464
    mem[3354] <= 16'h216f; // 0x80003468
    mem[3355] <= 16'h6e28; // 0x8000346c
    mem[3356] <= 16'h296c; // 0x80003470
    mem[3357] <= 16'h7325; // 0x80003474
    mem[3358] <= 16'h2520; // 0x80003478
    mem[3359] <= 16'h0000; // 0x8000347c
 
 
//================================================================
//== Section  .eh_frame
//================================================================
    mem[3360] <= 16'h0010; // 0x80003480
    mem[3361] <= 16'h0000; // 0x80003484
    mem[3362] <= 16'h7a03; // 0x80003488
    mem[3363] <= 16'h7c01; // 0x8000348c
    mem[3364] <= 16'h0c1b; // 0x80003490
    mem[3365] <= 16'h0010; // 0x80003494
    mem[3366] <= 16'h0018; // 0x80003498
    mem[3367] <= 16'hf2e8; // 0x8000349c
    mem[3368] <= 16'h0474; // 0x800034a0
    mem[3369] <= 16'h0000; // 0x800034a4
    mem[3370] <= 16'h0010; // 0x800034a8
    mem[3371] <= 16'h002c; // 0x800034ac
    mem[3372] <= 16'hf748; // 0x800034b0
    mem[3373] <= 16'h0428; // 0x800034b4
    mem[3374] <= 16'h0000; // 0x800034b8
 
 
end
endmodule
